module pe_top (state, rdpix, addrpix, valid, reset );
	input [1023:0] 	state;
	input        	rdpix;
	output [9:0] 	addrpix;
	output [1023:0] 	reset;
	output        	valid;
// Level 0
wire [1023:0] state_0;
wire [1023:0] reset_0;
wire [1023:0] ctrlreset_0;
wire [255:0] enable_0;
wire [255:0] rdpix_0;
wire [255:0] valid_0;
wire [511:0] addrpix_0;
	pe #(.ADR_WIDTH(2)) pe_0_0 (.state(state_0[3:0]),.ctrlreset(ctrlreset_0[3:0]),.reset(reset_0[3:0]),.enable(enable_0[0]),.valid(valid_0[0]),.rdpix(rdpix_0[0]),.addrpix({addrpix_0[256],addrpix_0[0]}));
	pe #(.ADR_WIDTH(2)) pe_0_1 (.state(state_0[7:4]),.ctrlreset(ctrlreset_0[7:4]),.reset(reset_0[7:4]),.enable(enable_0[1]),.valid(valid_0[1]),.rdpix(rdpix_0[1]),.addrpix({addrpix_0[257],addrpix_0[1]}));
	pe #(.ADR_WIDTH(2)) pe_0_2 (.state(state_0[11:8]),.ctrlreset(ctrlreset_0[11:8]),.reset(reset_0[11:8]),.enable(enable_0[2]),.valid(valid_0[2]),.rdpix(rdpix_0[2]),.addrpix({addrpix_0[258],addrpix_0[2]}));
	pe #(.ADR_WIDTH(2)) pe_0_3 (.state(state_0[15:12]),.ctrlreset(ctrlreset_0[15:12]),.reset(reset_0[15:12]),.enable(enable_0[3]),.valid(valid_0[3]),.rdpix(rdpix_0[3]),.addrpix({addrpix_0[259],addrpix_0[3]}));
	pe #(.ADR_WIDTH(2)) pe_0_4 (.state(state_0[19:16]),.ctrlreset(ctrlreset_0[19:16]),.reset(reset_0[19:16]),.enable(enable_0[4]),.valid(valid_0[4]),.rdpix(rdpix_0[4]),.addrpix({addrpix_0[260],addrpix_0[4]}));
	pe #(.ADR_WIDTH(2)) pe_0_5 (.state(state_0[23:20]),.ctrlreset(ctrlreset_0[23:20]),.reset(reset_0[23:20]),.enable(enable_0[5]),.valid(valid_0[5]),.rdpix(rdpix_0[5]),.addrpix({addrpix_0[261],addrpix_0[5]}));
	pe #(.ADR_WIDTH(2)) pe_0_6 (.state(state_0[27:24]),.ctrlreset(ctrlreset_0[27:24]),.reset(reset_0[27:24]),.enable(enable_0[6]),.valid(valid_0[6]),.rdpix(rdpix_0[6]),.addrpix({addrpix_0[262],addrpix_0[6]}));
	pe #(.ADR_WIDTH(2)) pe_0_7 (.state(state_0[31:28]),.ctrlreset(ctrlreset_0[31:28]),.reset(reset_0[31:28]),.enable(enable_0[7]),.valid(valid_0[7]),.rdpix(rdpix_0[7]),.addrpix({addrpix_0[263],addrpix_0[7]}));
	pe #(.ADR_WIDTH(2)) pe_0_8 (.state(state_0[35:32]),.ctrlreset(ctrlreset_0[35:32]),.reset(reset_0[35:32]),.enable(enable_0[8]),.valid(valid_0[8]),.rdpix(rdpix_0[8]),.addrpix({addrpix_0[264],addrpix_0[8]}));
	pe #(.ADR_WIDTH(2)) pe_0_9 (.state(state_0[39:36]),.ctrlreset(ctrlreset_0[39:36]),.reset(reset_0[39:36]),.enable(enable_0[9]),.valid(valid_0[9]),.rdpix(rdpix_0[9]),.addrpix({addrpix_0[265],addrpix_0[9]}));
	pe #(.ADR_WIDTH(2)) pe_0_10 (.state(state_0[43:40]),.ctrlreset(ctrlreset_0[43:40]),.reset(reset_0[43:40]),.enable(enable_0[10]),.valid(valid_0[10]),.rdpix(rdpix_0[10]),.addrpix({addrpix_0[266],addrpix_0[10]}));
	pe #(.ADR_WIDTH(2)) pe_0_11 (.state(state_0[47:44]),.ctrlreset(ctrlreset_0[47:44]),.reset(reset_0[47:44]),.enable(enable_0[11]),.valid(valid_0[11]),.rdpix(rdpix_0[11]),.addrpix({addrpix_0[267],addrpix_0[11]}));
	pe #(.ADR_WIDTH(2)) pe_0_12 (.state(state_0[51:48]),.ctrlreset(ctrlreset_0[51:48]),.reset(reset_0[51:48]),.enable(enable_0[12]),.valid(valid_0[12]),.rdpix(rdpix_0[12]),.addrpix({addrpix_0[268],addrpix_0[12]}));
	pe #(.ADR_WIDTH(2)) pe_0_13 (.state(state_0[55:52]),.ctrlreset(ctrlreset_0[55:52]),.reset(reset_0[55:52]),.enable(enable_0[13]),.valid(valid_0[13]),.rdpix(rdpix_0[13]),.addrpix({addrpix_0[269],addrpix_0[13]}));
	pe #(.ADR_WIDTH(2)) pe_0_14 (.state(state_0[59:56]),.ctrlreset(ctrlreset_0[59:56]),.reset(reset_0[59:56]),.enable(enable_0[14]),.valid(valid_0[14]),.rdpix(rdpix_0[14]),.addrpix({addrpix_0[270],addrpix_0[14]}));
	pe #(.ADR_WIDTH(2)) pe_0_15 (.state(state_0[63:60]),.ctrlreset(ctrlreset_0[63:60]),.reset(reset_0[63:60]),.enable(enable_0[15]),.valid(valid_0[15]),.rdpix(rdpix_0[15]),.addrpix({addrpix_0[271],addrpix_0[15]}));
	pe #(.ADR_WIDTH(2)) pe_0_16 (.state(state_0[67:64]),.ctrlreset(ctrlreset_0[67:64]),.reset(reset_0[67:64]),.enable(enable_0[16]),.valid(valid_0[16]),.rdpix(rdpix_0[16]),.addrpix({addrpix_0[272],addrpix_0[16]}));
	pe #(.ADR_WIDTH(2)) pe_0_17 (.state(state_0[71:68]),.ctrlreset(ctrlreset_0[71:68]),.reset(reset_0[71:68]),.enable(enable_0[17]),.valid(valid_0[17]),.rdpix(rdpix_0[17]),.addrpix({addrpix_0[273],addrpix_0[17]}));
	pe #(.ADR_WIDTH(2)) pe_0_18 (.state(state_0[75:72]),.ctrlreset(ctrlreset_0[75:72]),.reset(reset_0[75:72]),.enable(enable_0[18]),.valid(valid_0[18]),.rdpix(rdpix_0[18]),.addrpix({addrpix_0[274],addrpix_0[18]}));
	pe #(.ADR_WIDTH(2)) pe_0_19 (.state(state_0[79:76]),.ctrlreset(ctrlreset_0[79:76]),.reset(reset_0[79:76]),.enable(enable_0[19]),.valid(valid_0[19]),.rdpix(rdpix_0[19]),.addrpix({addrpix_0[275],addrpix_0[19]}));
	pe #(.ADR_WIDTH(2)) pe_0_20 (.state(state_0[83:80]),.ctrlreset(ctrlreset_0[83:80]),.reset(reset_0[83:80]),.enable(enable_0[20]),.valid(valid_0[20]),.rdpix(rdpix_0[20]),.addrpix({addrpix_0[276],addrpix_0[20]}));
	pe #(.ADR_WIDTH(2)) pe_0_21 (.state(state_0[87:84]),.ctrlreset(ctrlreset_0[87:84]),.reset(reset_0[87:84]),.enable(enable_0[21]),.valid(valid_0[21]),.rdpix(rdpix_0[21]),.addrpix({addrpix_0[277],addrpix_0[21]}));
	pe #(.ADR_WIDTH(2)) pe_0_22 (.state(state_0[91:88]),.ctrlreset(ctrlreset_0[91:88]),.reset(reset_0[91:88]),.enable(enable_0[22]),.valid(valid_0[22]),.rdpix(rdpix_0[22]),.addrpix({addrpix_0[278],addrpix_0[22]}));
	pe #(.ADR_WIDTH(2)) pe_0_23 (.state(state_0[95:92]),.ctrlreset(ctrlreset_0[95:92]),.reset(reset_0[95:92]),.enable(enable_0[23]),.valid(valid_0[23]),.rdpix(rdpix_0[23]),.addrpix({addrpix_0[279],addrpix_0[23]}));
	pe #(.ADR_WIDTH(2)) pe_0_24 (.state(state_0[99:96]),.ctrlreset(ctrlreset_0[99:96]),.reset(reset_0[99:96]),.enable(enable_0[24]),.valid(valid_0[24]),.rdpix(rdpix_0[24]),.addrpix({addrpix_0[280],addrpix_0[24]}));
	pe #(.ADR_WIDTH(2)) pe_0_25 (.state(state_0[103:100]),.ctrlreset(ctrlreset_0[103:100]),.reset(reset_0[103:100]),.enable(enable_0[25]),.valid(valid_0[25]),.rdpix(rdpix_0[25]),.addrpix({addrpix_0[281],addrpix_0[25]}));
	pe #(.ADR_WIDTH(2)) pe_0_26 (.state(state_0[107:104]),.ctrlreset(ctrlreset_0[107:104]),.reset(reset_0[107:104]),.enable(enable_0[26]),.valid(valid_0[26]),.rdpix(rdpix_0[26]),.addrpix({addrpix_0[282],addrpix_0[26]}));
	pe #(.ADR_WIDTH(2)) pe_0_27 (.state(state_0[111:108]),.ctrlreset(ctrlreset_0[111:108]),.reset(reset_0[111:108]),.enable(enable_0[27]),.valid(valid_0[27]),.rdpix(rdpix_0[27]),.addrpix({addrpix_0[283],addrpix_0[27]}));
	pe #(.ADR_WIDTH(2)) pe_0_28 (.state(state_0[115:112]),.ctrlreset(ctrlreset_0[115:112]),.reset(reset_0[115:112]),.enable(enable_0[28]),.valid(valid_0[28]),.rdpix(rdpix_0[28]),.addrpix({addrpix_0[284],addrpix_0[28]}));
	pe #(.ADR_WIDTH(2)) pe_0_29 (.state(state_0[119:116]),.ctrlreset(ctrlreset_0[119:116]),.reset(reset_0[119:116]),.enable(enable_0[29]),.valid(valid_0[29]),.rdpix(rdpix_0[29]),.addrpix({addrpix_0[285],addrpix_0[29]}));
	pe #(.ADR_WIDTH(2)) pe_0_30 (.state(state_0[123:120]),.ctrlreset(ctrlreset_0[123:120]),.reset(reset_0[123:120]),.enable(enable_0[30]),.valid(valid_0[30]),.rdpix(rdpix_0[30]),.addrpix({addrpix_0[286],addrpix_0[30]}));
	pe #(.ADR_WIDTH(2)) pe_0_31 (.state(state_0[127:124]),.ctrlreset(ctrlreset_0[127:124]),.reset(reset_0[127:124]),.enable(enable_0[31]),.valid(valid_0[31]),.rdpix(rdpix_0[31]),.addrpix({addrpix_0[287],addrpix_0[31]}));
	pe #(.ADR_WIDTH(2)) pe_0_32 (.state(state_0[131:128]),.ctrlreset(ctrlreset_0[131:128]),.reset(reset_0[131:128]),.enable(enable_0[32]),.valid(valid_0[32]),.rdpix(rdpix_0[32]),.addrpix({addrpix_0[288],addrpix_0[32]}));
	pe #(.ADR_WIDTH(2)) pe_0_33 (.state(state_0[135:132]),.ctrlreset(ctrlreset_0[135:132]),.reset(reset_0[135:132]),.enable(enable_0[33]),.valid(valid_0[33]),.rdpix(rdpix_0[33]),.addrpix({addrpix_0[289],addrpix_0[33]}));
	pe #(.ADR_WIDTH(2)) pe_0_34 (.state(state_0[139:136]),.ctrlreset(ctrlreset_0[139:136]),.reset(reset_0[139:136]),.enable(enable_0[34]),.valid(valid_0[34]),.rdpix(rdpix_0[34]),.addrpix({addrpix_0[290],addrpix_0[34]}));
	pe #(.ADR_WIDTH(2)) pe_0_35 (.state(state_0[143:140]),.ctrlreset(ctrlreset_0[143:140]),.reset(reset_0[143:140]),.enable(enable_0[35]),.valid(valid_0[35]),.rdpix(rdpix_0[35]),.addrpix({addrpix_0[291],addrpix_0[35]}));
	pe #(.ADR_WIDTH(2)) pe_0_36 (.state(state_0[147:144]),.ctrlreset(ctrlreset_0[147:144]),.reset(reset_0[147:144]),.enable(enable_0[36]),.valid(valid_0[36]),.rdpix(rdpix_0[36]),.addrpix({addrpix_0[292],addrpix_0[36]}));
	pe #(.ADR_WIDTH(2)) pe_0_37 (.state(state_0[151:148]),.ctrlreset(ctrlreset_0[151:148]),.reset(reset_0[151:148]),.enable(enable_0[37]),.valid(valid_0[37]),.rdpix(rdpix_0[37]),.addrpix({addrpix_0[293],addrpix_0[37]}));
	pe #(.ADR_WIDTH(2)) pe_0_38 (.state(state_0[155:152]),.ctrlreset(ctrlreset_0[155:152]),.reset(reset_0[155:152]),.enable(enable_0[38]),.valid(valid_0[38]),.rdpix(rdpix_0[38]),.addrpix({addrpix_0[294],addrpix_0[38]}));
	pe #(.ADR_WIDTH(2)) pe_0_39 (.state(state_0[159:156]),.ctrlreset(ctrlreset_0[159:156]),.reset(reset_0[159:156]),.enable(enable_0[39]),.valid(valid_0[39]),.rdpix(rdpix_0[39]),.addrpix({addrpix_0[295],addrpix_0[39]}));
	pe #(.ADR_WIDTH(2)) pe_0_40 (.state(state_0[163:160]),.ctrlreset(ctrlreset_0[163:160]),.reset(reset_0[163:160]),.enable(enable_0[40]),.valid(valid_0[40]),.rdpix(rdpix_0[40]),.addrpix({addrpix_0[296],addrpix_0[40]}));
	pe #(.ADR_WIDTH(2)) pe_0_41 (.state(state_0[167:164]),.ctrlreset(ctrlreset_0[167:164]),.reset(reset_0[167:164]),.enable(enable_0[41]),.valid(valid_0[41]),.rdpix(rdpix_0[41]),.addrpix({addrpix_0[297],addrpix_0[41]}));
	pe #(.ADR_WIDTH(2)) pe_0_42 (.state(state_0[171:168]),.ctrlreset(ctrlreset_0[171:168]),.reset(reset_0[171:168]),.enable(enable_0[42]),.valid(valid_0[42]),.rdpix(rdpix_0[42]),.addrpix({addrpix_0[298],addrpix_0[42]}));
	pe #(.ADR_WIDTH(2)) pe_0_43 (.state(state_0[175:172]),.ctrlreset(ctrlreset_0[175:172]),.reset(reset_0[175:172]),.enable(enable_0[43]),.valid(valid_0[43]),.rdpix(rdpix_0[43]),.addrpix({addrpix_0[299],addrpix_0[43]}));
	pe #(.ADR_WIDTH(2)) pe_0_44 (.state(state_0[179:176]),.ctrlreset(ctrlreset_0[179:176]),.reset(reset_0[179:176]),.enable(enable_0[44]),.valid(valid_0[44]),.rdpix(rdpix_0[44]),.addrpix({addrpix_0[300],addrpix_0[44]}));
	pe #(.ADR_WIDTH(2)) pe_0_45 (.state(state_0[183:180]),.ctrlreset(ctrlreset_0[183:180]),.reset(reset_0[183:180]),.enable(enable_0[45]),.valid(valid_0[45]),.rdpix(rdpix_0[45]),.addrpix({addrpix_0[301],addrpix_0[45]}));
	pe #(.ADR_WIDTH(2)) pe_0_46 (.state(state_0[187:184]),.ctrlreset(ctrlreset_0[187:184]),.reset(reset_0[187:184]),.enable(enable_0[46]),.valid(valid_0[46]),.rdpix(rdpix_0[46]),.addrpix({addrpix_0[302],addrpix_0[46]}));
	pe #(.ADR_WIDTH(2)) pe_0_47 (.state(state_0[191:188]),.ctrlreset(ctrlreset_0[191:188]),.reset(reset_0[191:188]),.enable(enable_0[47]),.valid(valid_0[47]),.rdpix(rdpix_0[47]),.addrpix({addrpix_0[303],addrpix_0[47]}));
	pe #(.ADR_WIDTH(2)) pe_0_48 (.state(state_0[195:192]),.ctrlreset(ctrlreset_0[195:192]),.reset(reset_0[195:192]),.enable(enable_0[48]),.valid(valid_0[48]),.rdpix(rdpix_0[48]),.addrpix({addrpix_0[304],addrpix_0[48]}));
	pe #(.ADR_WIDTH(2)) pe_0_49 (.state(state_0[199:196]),.ctrlreset(ctrlreset_0[199:196]),.reset(reset_0[199:196]),.enable(enable_0[49]),.valid(valid_0[49]),.rdpix(rdpix_0[49]),.addrpix({addrpix_0[305],addrpix_0[49]}));
	pe #(.ADR_WIDTH(2)) pe_0_50 (.state(state_0[203:200]),.ctrlreset(ctrlreset_0[203:200]),.reset(reset_0[203:200]),.enable(enable_0[50]),.valid(valid_0[50]),.rdpix(rdpix_0[50]),.addrpix({addrpix_0[306],addrpix_0[50]}));
	pe #(.ADR_WIDTH(2)) pe_0_51 (.state(state_0[207:204]),.ctrlreset(ctrlreset_0[207:204]),.reset(reset_0[207:204]),.enable(enable_0[51]),.valid(valid_0[51]),.rdpix(rdpix_0[51]),.addrpix({addrpix_0[307],addrpix_0[51]}));
	pe #(.ADR_WIDTH(2)) pe_0_52 (.state(state_0[211:208]),.ctrlreset(ctrlreset_0[211:208]),.reset(reset_0[211:208]),.enable(enable_0[52]),.valid(valid_0[52]),.rdpix(rdpix_0[52]),.addrpix({addrpix_0[308],addrpix_0[52]}));
	pe #(.ADR_WIDTH(2)) pe_0_53 (.state(state_0[215:212]),.ctrlreset(ctrlreset_0[215:212]),.reset(reset_0[215:212]),.enable(enable_0[53]),.valid(valid_0[53]),.rdpix(rdpix_0[53]),.addrpix({addrpix_0[309],addrpix_0[53]}));
	pe #(.ADR_WIDTH(2)) pe_0_54 (.state(state_0[219:216]),.ctrlreset(ctrlreset_0[219:216]),.reset(reset_0[219:216]),.enable(enable_0[54]),.valid(valid_0[54]),.rdpix(rdpix_0[54]),.addrpix({addrpix_0[310],addrpix_0[54]}));
	pe #(.ADR_WIDTH(2)) pe_0_55 (.state(state_0[223:220]),.ctrlreset(ctrlreset_0[223:220]),.reset(reset_0[223:220]),.enable(enable_0[55]),.valid(valid_0[55]),.rdpix(rdpix_0[55]),.addrpix({addrpix_0[311],addrpix_0[55]}));
	pe #(.ADR_WIDTH(2)) pe_0_56 (.state(state_0[227:224]),.ctrlreset(ctrlreset_0[227:224]),.reset(reset_0[227:224]),.enable(enable_0[56]),.valid(valid_0[56]),.rdpix(rdpix_0[56]),.addrpix({addrpix_0[312],addrpix_0[56]}));
	pe #(.ADR_WIDTH(2)) pe_0_57 (.state(state_0[231:228]),.ctrlreset(ctrlreset_0[231:228]),.reset(reset_0[231:228]),.enable(enable_0[57]),.valid(valid_0[57]),.rdpix(rdpix_0[57]),.addrpix({addrpix_0[313],addrpix_0[57]}));
	pe #(.ADR_WIDTH(2)) pe_0_58 (.state(state_0[235:232]),.ctrlreset(ctrlreset_0[235:232]),.reset(reset_0[235:232]),.enable(enable_0[58]),.valid(valid_0[58]),.rdpix(rdpix_0[58]),.addrpix({addrpix_0[314],addrpix_0[58]}));
	pe #(.ADR_WIDTH(2)) pe_0_59 (.state(state_0[239:236]),.ctrlreset(ctrlreset_0[239:236]),.reset(reset_0[239:236]),.enable(enable_0[59]),.valid(valid_0[59]),.rdpix(rdpix_0[59]),.addrpix({addrpix_0[315],addrpix_0[59]}));
	pe #(.ADR_WIDTH(2)) pe_0_60 (.state(state_0[243:240]),.ctrlreset(ctrlreset_0[243:240]),.reset(reset_0[243:240]),.enable(enable_0[60]),.valid(valid_0[60]),.rdpix(rdpix_0[60]),.addrpix({addrpix_0[316],addrpix_0[60]}));
	pe #(.ADR_WIDTH(2)) pe_0_61 (.state(state_0[247:244]),.ctrlreset(ctrlreset_0[247:244]),.reset(reset_0[247:244]),.enable(enable_0[61]),.valid(valid_0[61]),.rdpix(rdpix_0[61]),.addrpix({addrpix_0[317],addrpix_0[61]}));
	pe #(.ADR_WIDTH(2)) pe_0_62 (.state(state_0[251:248]),.ctrlreset(ctrlreset_0[251:248]),.reset(reset_0[251:248]),.enable(enable_0[62]),.valid(valid_0[62]),.rdpix(rdpix_0[62]),.addrpix({addrpix_0[318],addrpix_0[62]}));
	pe #(.ADR_WIDTH(2)) pe_0_63 (.state(state_0[255:252]),.ctrlreset(ctrlreset_0[255:252]),.reset(reset_0[255:252]),.enable(enable_0[63]),.valid(valid_0[63]),.rdpix(rdpix_0[63]),.addrpix({addrpix_0[319],addrpix_0[63]}));
	pe #(.ADR_WIDTH(2)) pe_0_64 (.state(state_0[259:256]),.ctrlreset(ctrlreset_0[259:256]),.reset(reset_0[259:256]),.enable(enable_0[64]),.valid(valid_0[64]),.rdpix(rdpix_0[64]),.addrpix({addrpix_0[320],addrpix_0[64]}));
	pe #(.ADR_WIDTH(2)) pe_0_65 (.state(state_0[263:260]),.ctrlreset(ctrlreset_0[263:260]),.reset(reset_0[263:260]),.enable(enable_0[65]),.valid(valid_0[65]),.rdpix(rdpix_0[65]),.addrpix({addrpix_0[321],addrpix_0[65]}));
	pe #(.ADR_WIDTH(2)) pe_0_66 (.state(state_0[267:264]),.ctrlreset(ctrlreset_0[267:264]),.reset(reset_0[267:264]),.enable(enable_0[66]),.valid(valid_0[66]),.rdpix(rdpix_0[66]),.addrpix({addrpix_0[322],addrpix_0[66]}));
	pe #(.ADR_WIDTH(2)) pe_0_67 (.state(state_0[271:268]),.ctrlreset(ctrlreset_0[271:268]),.reset(reset_0[271:268]),.enable(enable_0[67]),.valid(valid_0[67]),.rdpix(rdpix_0[67]),.addrpix({addrpix_0[323],addrpix_0[67]}));
	pe #(.ADR_WIDTH(2)) pe_0_68 (.state(state_0[275:272]),.ctrlreset(ctrlreset_0[275:272]),.reset(reset_0[275:272]),.enable(enable_0[68]),.valid(valid_0[68]),.rdpix(rdpix_0[68]),.addrpix({addrpix_0[324],addrpix_0[68]}));
	pe #(.ADR_WIDTH(2)) pe_0_69 (.state(state_0[279:276]),.ctrlreset(ctrlreset_0[279:276]),.reset(reset_0[279:276]),.enable(enable_0[69]),.valid(valid_0[69]),.rdpix(rdpix_0[69]),.addrpix({addrpix_0[325],addrpix_0[69]}));
	pe #(.ADR_WIDTH(2)) pe_0_70 (.state(state_0[283:280]),.ctrlreset(ctrlreset_0[283:280]),.reset(reset_0[283:280]),.enable(enable_0[70]),.valid(valid_0[70]),.rdpix(rdpix_0[70]),.addrpix({addrpix_0[326],addrpix_0[70]}));
	pe #(.ADR_WIDTH(2)) pe_0_71 (.state(state_0[287:284]),.ctrlreset(ctrlreset_0[287:284]),.reset(reset_0[287:284]),.enable(enable_0[71]),.valid(valid_0[71]),.rdpix(rdpix_0[71]),.addrpix({addrpix_0[327],addrpix_0[71]}));
	pe #(.ADR_WIDTH(2)) pe_0_72 (.state(state_0[291:288]),.ctrlreset(ctrlreset_0[291:288]),.reset(reset_0[291:288]),.enable(enable_0[72]),.valid(valid_0[72]),.rdpix(rdpix_0[72]),.addrpix({addrpix_0[328],addrpix_0[72]}));
	pe #(.ADR_WIDTH(2)) pe_0_73 (.state(state_0[295:292]),.ctrlreset(ctrlreset_0[295:292]),.reset(reset_0[295:292]),.enable(enable_0[73]),.valid(valid_0[73]),.rdpix(rdpix_0[73]),.addrpix({addrpix_0[329],addrpix_0[73]}));
	pe #(.ADR_WIDTH(2)) pe_0_74 (.state(state_0[299:296]),.ctrlreset(ctrlreset_0[299:296]),.reset(reset_0[299:296]),.enable(enable_0[74]),.valid(valid_0[74]),.rdpix(rdpix_0[74]),.addrpix({addrpix_0[330],addrpix_0[74]}));
	pe #(.ADR_WIDTH(2)) pe_0_75 (.state(state_0[303:300]),.ctrlreset(ctrlreset_0[303:300]),.reset(reset_0[303:300]),.enable(enable_0[75]),.valid(valid_0[75]),.rdpix(rdpix_0[75]),.addrpix({addrpix_0[331],addrpix_0[75]}));
	pe #(.ADR_WIDTH(2)) pe_0_76 (.state(state_0[307:304]),.ctrlreset(ctrlreset_0[307:304]),.reset(reset_0[307:304]),.enable(enable_0[76]),.valid(valid_0[76]),.rdpix(rdpix_0[76]),.addrpix({addrpix_0[332],addrpix_0[76]}));
	pe #(.ADR_WIDTH(2)) pe_0_77 (.state(state_0[311:308]),.ctrlreset(ctrlreset_0[311:308]),.reset(reset_0[311:308]),.enable(enable_0[77]),.valid(valid_0[77]),.rdpix(rdpix_0[77]),.addrpix({addrpix_0[333],addrpix_0[77]}));
	pe #(.ADR_WIDTH(2)) pe_0_78 (.state(state_0[315:312]),.ctrlreset(ctrlreset_0[315:312]),.reset(reset_0[315:312]),.enable(enable_0[78]),.valid(valid_0[78]),.rdpix(rdpix_0[78]),.addrpix({addrpix_0[334],addrpix_0[78]}));
	pe #(.ADR_WIDTH(2)) pe_0_79 (.state(state_0[319:316]),.ctrlreset(ctrlreset_0[319:316]),.reset(reset_0[319:316]),.enable(enable_0[79]),.valid(valid_0[79]),.rdpix(rdpix_0[79]),.addrpix({addrpix_0[335],addrpix_0[79]}));
	pe #(.ADR_WIDTH(2)) pe_0_80 (.state(state_0[323:320]),.ctrlreset(ctrlreset_0[323:320]),.reset(reset_0[323:320]),.enable(enable_0[80]),.valid(valid_0[80]),.rdpix(rdpix_0[80]),.addrpix({addrpix_0[336],addrpix_0[80]}));
	pe #(.ADR_WIDTH(2)) pe_0_81 (.state(state_0[327:324]),.ctrlreset(ctrlreset_0[327:324]),.reset(reset_0[327:324]),.enable(enable_0[81]),.valid(valid_0[81]),.rdpix(rdpix_0[81]),.addrpix({addrpix_0[337],addrpix_0[81]}));
	pe #(.ADR_WIDTH(2)) pe_0_82 (.state(state_0[331:328]),.ctrlreset(ctrlreset_0[331:328]),.reset(reset_0[331:328]),.enable(enable_0[82]),.valid(valid_0[82]),.rdpix(rdpix_0[82]),.addrpix({addrpix_0[338],addrpix_0[82]}));
	pe #(.ADR_WIDTH(2)) pe_0_83 (.state(state_0[335:332]),.ctrlreset(ctrlreset_0[335:332]),.reset(reset_0[335:332]),.enable(enable_0[83]),.valid(valid_0[83]),.rdpix(rdpix_0[83]),.addrpix({addrpix_0[339],addrpix_0[83]}));
	pe #(.ADR_WIDTH(2)) pe_0_84 (.state(state_0[339:336]),.ctrlreset(ctrlreset_0[339:336]),.reset(reset_0[339:336]),.enable(enable_0[84]),.valid(valid_0[84]),.rdpix(rdpix_0[84]),.addrpix({addrpix_0[340],addrpix_0[84]}));
	pe #(.ADR_WIDTH(2)) pe_0_85 (.state(state_0[343:340]),.ctrlreset(ctrlreset_0[343:340]),.reset(reset_0[343:340]),.enable(enable_0[85]),.valid(valid_0[85]),.rdpix(rdpix_0[85]),.addrpix({addrpix_0[341],addrpix_0[85]}));
	pe #(.ADR_WIDTH(2)) pe_0_86 (.state(state_0[347:344]),.ctrlreset(ctrlreset_0[347:344]),.reset(reset_0[347:344]),.enable(enable_0[86]),.valid(valid_0[86]),.rdpix(rdpix_0[86]),.addrpix({addrpix_0[342],addrpix_0[86]}));
	pe #(.ADR_WIDTH(2)) pe_0_87 (.state(state_0[351:348]),.ctrlreset(ctrlreset_0[351:348]),.reset(reset_0[351:348]),.enable(enable_0[87]),.valid(valid_0[87]),.rdpix(rdpix_0[87]),.addrpix({addrpix_0[343],addrpix_0[87]}));
	pe #(.ADR_WIDTH(2)) pe_0_88 (.state(state_0[355:352]),.ctrlreset(ctrlreset_0[355:352]),.reset(reset_0[355:352]),.enable(enable_0[88]),.valid(valid_0[88]),.rdpix(rdpix_0[88]),.addrpix({addrpix_0[344],addrpix_0[88]}));
	pe #(.ADR_WIDTH(2)) pe_0_89 (.state(state_0[359:356]),.ctrlreset(ctrlreset_0[359:356]),.reset(reset_0[359:356]),.enable(enable_0[89]),.valid(valid_0[89]),.rdpix(rdpix_0[89]),.addrpix({addrpix_0[345],addrpix_0[89]}));
	pe #(.ADR_WIDTH(2)) pe_0_90 (.state(state_0[363:360]),.ctrlreset(ctrlreset_0[363:360]),.reset(reset_0[363:360]),.enable(enable_0[90]),.valid(valid_0[90]),.rdpix(rdpix_0[90]),.addrpix({addrpix_0[346],addrpix_0[90]}));
	pe #(.ADR_WIDTH(2)) pe_0_91 (.state(state_0[367:364]),.ctrlreset(ctrlreset_0[367:364]),.reset(reset_0[367:364]),.enable(enable_0[91]),.valid(valid_0[91]),.rdpix(rdpix_0[91]),.addrpix({addrpix_0[347],addrpix_0[91]}));
	pe #(.ADR_WIDTH(2)) pe_0_92 (.state(state_0[371:368]),.ctrlreset(ctrlreset_0[371:368]),.reset(reset_0[371:368]),.enable(enable_0[92]),.valid(valid_0[92]),.rdpix(rdpix_0[92]),.addrpix({addrpix_0[348],addrpix_0[92]}));
	pe #(.ADR_WIDTH(2)) pe_0_93 (.state(state_0[375:372]),.ctrlreset(ctrlreset_0[375:372]),.reset(reset_0[375:372]),.enable(enable_0[93]),.valid(valid_0[93]),.rdpix(rdpix_0[93]),.addrpix({addrpix_0[349],addrpix_0[93]}));
	pe #(.ADR_WIDTH(2)) pe_0_94 (.state(state_0[379:376]),.ctrlreset(ctrlreset_0[379:376]),.reset(reset_0[379:376]),.enable(enable_0[94]),.valid(valid_0[94]),.rdpix(rdpix_0[94]),.addrpix({addrpix_0[350],addrpix_0[94]}));
	pe #(.ADR_WIDTH(2)) pe_0_95 (.state(state_0[383:380]),.ctrlreset(ctrlreset_0[383:380]),.reset(reset_0[383:380]),.enable(enable_0[95]),.valid(valid_0[95]),.rdpix(rdpix_0[95]),.addrpix({addrpix_0[351],addrpix_0[95]}));
	pe #(.ADR_WIDTH(2)) pe_0_96 (.state(state_0[387:384]),.ctrlreset(ctrlreset_0[387:384]),.reset(reset_0[387:384]),.enable(enable_0[96]),.valid(valid_0[96]),.rdpix(rdpix_0[96]),.addrpix({addrpix_0[352],addrpix_0[96]}));
	pe #(.ADR_WIDTH(2)) pe_0_97 (.state(state_0[391:388]),.ctrlreset(ctrlreset_0[391:388]),.reset(reset_0[391:388]),.enable(enable_0[97]),.valid(valid_0[97]),.rdpix(rdpix_0[97]),.addrpix({addrpix_0[353],addrpix_0[97]}));
	pe #(.ADR_WIDTH(2)) pe_0_98 (.state(state_0[395:392]),.ctrlreset(ctrlreset_0[395:392]),.reset(reset_0[395:392]),.enable(enable_0[98]),.valid(valid_0[98]),.rdpix(rdpix_0[98]),.addrpix({addrpix_0[354],addrpix_0[98]}));
	pe #(.ADR_WIDTH(2)) pe_0_99 (.state(state_0[399:396]),.ctrlreset(ctrlreset_0[399:396]),.reset(reset_0[399:396]),.enable(enable_0[99]),.valid(valid_0[99]),.rdpix(rdpix_0[99]),.addrpix({addrpix_0[355],addrpix_0[99]}));
	pe #(.ADR_WIDTH(2)) pe_0_100 (.state(state_0[403:400]),.ctrlreset(ctrlreset_0[403:400]),.reset(reset_0[403:400]),.enable(enable_0[100]),.valid(valid_0[100]),.rdpix(rdpix_0[100]),.addrpix({addrpix_0[356],addrpix_0[100]}));
	pe #(.ADR_WIDTH(2)) pe_0_101 (.state(state_0[407:404]),.ctrlreset(ctrlreset_0[407:404]),.reset(reset_0[407:404]),.enable(enable_0[101]),.valid(valid_0[101]),.rdpix(rdpix_0[101]),.addrpix({addrpix_0[357],addrpix_0[101]}));
	pe #(.ADR_WIDTH(2)) pe_0_102 (.state(state_0[411:408]),.ctrlreset(ctrlreset_0[411:408]),.reset(reset_0[411:408]),.enable(enable_0[102]),.valid(valid_0[102]),.rdpix(rdpix_0[102]),.addrpix({addrpix_0[358],addrpix_0[102]}));
	pe #(.ADR_WIDTH(2)) pe_0_103 (.state(state_0[415:412]),.ctrlreset(ctrlreset_0[415:412]),.reset(reset_0[415:412]),.enable(enable_0[103]),.valid(valid_0[103]),.rdpix(rdpix_0[103]),.addrpix({addrpix_0[359],addrpix_0[103]}));
	pe #(.ADR_WIDTH(2)) pe_0_104 (.state(state_0[419:416]),.ctrlreset(ctrlreset_0[419:416]),.reset(reset_0[419:416]),.enable(enable_0[104]),.valid(valid_0[104]),.rdpix(rdpix_0[104]),.addrpix({addrpix_0[360],addrpix_0[104]}));
	pe #(.ADR_WIDTH(2)) pe_0_105 (.state(state_0[423:420]),.ctrlreset(ctrlreset_0[423:420]),.reset(reset_0[423:420]),.enable(enable_0[105]),.valid(valid_0[105]),.rdpix(rdpix_0[105]),.addrpix({addrpix_0[361],addrpix_0[105]}));
	pe #(.ADR_WIDTH(2)) pe_0_106 (.state(state_0[427:424]),.ctrlreset(ctrlreset_0[427:424]),.reset(reset_0[427:424]),.enable(enable_0[106]),.valid(valid_0[106]),.rdpix(rdpix_0[106]),.addrpix({addrpix_0[362],addrpix_0[106]}));
	pe #(.ADR_WIDTH(2)) pe_0_107 (.state(state_0[431:428]),.ctrlreset(ctrlreset_0[431:428]),.reset(reset_0[431:428]),.enable(enable_0[107]),.valid(valid_0[107]),.rdpix(rdpix_0[107]),.addrpix({addrpix_0[363],addrpix_0[107]}));
	pe #(.ADR_WIDTH(2)) pe_0_108 (.state(state_0[435:432]),.ctrlreset(ctrlreset_0[435:432]),.reset(reset_0[435:432]),.enable(enable_0[108]),.valid(valid_0[108]),.rdpix(rdpix_0[108]),.addrpix({addrpix_0[364],addrpix_0[108]}));
	pe #(.ADR_WIDTH(2)) pe_0_109 (.state(state_0[439:436]),.ctrlreset(ctrlreset_0[439:436]),.reset(reset_0[439:436]),.enable(enable_0[109]),.valid(valid_0[109]),.rdpix(rdpix_0[109]),.addrpix({addrpix_0[365],addrpix_0[109]}));
	pe #(.ADR_WIDTH(2)) pe_0_110 (.state(state_0[443:440]),.ctrlreset(ctrlreset_0[443:440]),.reset(reset_0[443:440]),.enable(enable_0[110]),.valid(valid_0[110]),.rdpix(rdpix_0[110]),.addrpix({addrpix_0[366],addrpix_0[110]}));
	pe #(.ADR_WIDTH(2)) pe_0_111 (.state(state_0[447:444]),.ctrlreset(ctrlreset_0[447:444]),.reset(reset_0[447:444]),.enable(enable_0[111]),.valid(valid_0[111]),.rdpix(rdpix_0[111]),.addrpix({addrpix_0[367],addrpix_0[111]}));
	pe #(.ADR_WIDTH(2)) pe_0_112 (.state(state_0[451:448]),.ctrlreset(ctrlreset_0[451:448]),.reset(reset_0[451:448]),.enable(enable_0[112]),.valid(valid_0[112]),.rdpix(rdpix_0[112]),.addrpix({addrpix_0[368],addrpix_0[112]}));
	pe #(.ADR_WIDTH(2)) pe_0_113 (.state(state_0[455:452]),.ctrlreset(ctrlreset_0[455:452]),.reset(reset_0[455:452]),.enable(enable_0[113]),.valid(valid_0[113]),.rdpix(rdpix_0[113]),.addrpix({addrpix_0[369],addrpix_0[113]}));
	pe #(.ADR_WIDTH(2)) pe_0_114 (.state(state_0[459:456]),.ctrlreset(ctrlreset_0[459:456]),.reset(reset_0[459:456]),.enable(enable_0[114]),.valid(valid_0[114]),.rdpix(rdpix_0[114]),.addrpix({addrpix_0[370],addrpix_0[114]}));
	pe #(.ADR_WIDTH(2)) pe_0_115 (.state(state_0[463:460]),.ctrlreset(ctrlreset_0[463:460]),.reset(reset_0[463:460]),.enable(enable_0[115]),.valid(valid_0[115]),.rdpix(rdpix_0[115]),.addrpix({addrpix_0[371],addrpix_0[115]}));
	pe #(.ADR_WIDTH(2)) pe_0_116 (.state(state_0[467:464]),.ctrlreset(ctrlreset_0[467:464]),.reset(reset_0[467:464]),.enable(enable_0[116]),.valid(valid_0[116]),.rdpix(rdpix_0[116]),.addrpix({addrpix_0[372],addrpix_0[116]}));
	pe #(.ADR_WIDTH(2)) pe_0_117 (.state(state_0[471:468]),.ctrlreset(ctrlreset_0[471:468]),.reset(reset_0[471:468]),.enable(enable_0[117]),.valid(valid_0[117]),.rdpix(rdpix_0[117]),.addrpix({addrpix_0[373],addrpix_0[117]}));
	pe #(.ADR_WIDTH(2)) pe_0_118 (.state(state_0[475:472]),.ctrlreset(ctrlreset_0[475:472]),.reset(reset_0[475:472]),.enable(enable_0[118]),.valid(valid_0[118]),.rdpix(rdpix_0[118]),.addrpix({addrpix_0[374],addrpix_0[118]}));
	pe #(.ADR_WIDTH(2)) pe_0_119 (.state(state_0[479:476]),.ctrlreset(ctrlreset_0[479:476]),.reset(reset_0[479:476]),.enable(enable_0[119]),.valid(valid_0[119]),.rdpix(rdpix_0[119]),.addrpix({addrpix_0[375],addrpix_0[119]}));
	pe #(.ADR_WIDTH(2)) pe_0_120 (.state(state_0[483:480]),.ctrlreset(ctrlreset_0[483:480]),.reset(reset_0[483:480]),.enable(enable_0[120]),.valid(valid_0[120]),.rdpix(rdpix_0[120]),.addrpix({addrpix_0[376],addrpix_0[120]}));
	pe #(.ADR_WIDTH(2)) pe_0_121 (.state(state_0[487:484]),.ctrlreset(ctrlreset_0[487:484]),.reset(reset_0[487:484]),.enable(enable_0[121]),.valid(valid_0[121]),.rdpix(rdpix_0[121]),.addrpix({addrpix_0[377],addrpix_0[121]}));
	pe #(.ADR_WIDTH(2)) pe_0_122 (.state(state_0[491:488]),.ctrlreset(ctrlreset_0[491:488]),.reset(reset_0[491:488]),.enable(enable_0[122]),.valid(valid_0[122]),.rdpix(rdpix_0[122]),.addrpix({addrpix_0[378],addrpix_0[122]}));
	pe #(.ADR_WIDTH(2)) pe_0_123 (.state(state_0[495:492]),.ctrlreset(ctrlreset_0[495:492]),.reset(reset_0[495:492]),.enable(enable_0[123]),.valid(valid_0[123]),.rdpix(rdpix_0[123]),.addrpix({addrpix_0[379],addrpix_0[123]}));
	pe #(.ADR_WIDTH(2)) pe_0_124 (.state(state_0[499:496]),.ctrlreset(ctrlreset_0[499:496]),.reset(reset_0[499:496]),.enable(enable_0[124]),.valid(valid_0[124]),.rdpix(rdpix_0[124]),.addrpix({addrpix_0[380],addrpix_0[124]}));
	pe #(.ADR_WIDTH(2)) pe_0_125 (.state(state_0[503:500]),.ctrlreset(ctrlreset_0[503:500]),.reset(reset_0[503:500]),.enable(enable_0[125]),.valid(valid_0[125]),.rdpix(rdpix_0[125]),.addrpix({addrpix_0[381],addrpix_0[125]}));
	pe #(.ADR_WIDTH(2)) pe_0_126 (.state(state_0[507:504]),.ctrlreset(ctrlreset_0[507:504]),.reset(reset_0[507:504]),.enable(enable_0[126]),.valid(valid_0[126]),.rdpix(rdpix_0[126]),.addrpix({addrpix_0[382],addrpix_0[126]}));
	pe #(.ADR_WIDTH(2)) pe_0_127 (.state(state_0[511:508]),.ctrlreset(ctrlreset_0[511:508]),.reset(reset_0[511:508]),.enable(enable_0[127]),.valid(valid_0[127]),.rdpix(rdpix_0[127]),.addrpix({addrpix_0[383],addrpix_0[127]}));
	pe #(.ADR_WIDTH(2)) pe_0_128 (.state(state_0[515:512]),.ctrlreset(ctrlreset_0[515:512]),.reset(reset_0[515:512]),.enable(enable_0[128]),.valid(valid_0[128]),.rdpix(rdpix_0[128]),.addrpix({addrpix_0[384],addrpix_0[128]}));
	pe #(.ADR_WIDTH(2)) pe_0_129 (.state(state_0[519:516]),.ctrlreset(ctrlreset_0[519:516]),.reset(reset_0[519:516]),.enable(enable_0[129]),.valid(valid_0[129]),.rdpix(rdpix_0[129]),.addrpix({addrpix_0[385],addrpix_0[129]}));
	pe #(.ADR_WIDTH(2)) pe_0_130 (.state(state_0[523:520]),.ctrlreset(ctrlreset_0[523:520]),.reset(reset_0[523:520]),.enable(enable_0[130]),.valid(valid_0[130]),.rdpix(rdpix_0[130]),.addrpix({addrpix_0[386],addrpix_0[130]}));
	pe #(.ADR_WIDTH(2)) pe_0_131 (.state(state_0[527:524]),.ctrlreset(ctrlreset_0[527:524]),.reset(reset_0[527:524]),.enable(enable_0[131]),.valid(valid_0[131]),.rdpix(rdpix_0[131]),.addrpix({addrpix_0[387],addrpix_0[131]}));
	pe #(.ADR_WIDTH(2)) pe_0_132 (.state(state_0[531:528]),.ctrlreset(ctrlreset_0[531:528]),.reset(reset_0[531:528]),.enable(enable_0[132]),.valid(valid_0[132]),.rdpix(rdpix_0[132]),.addrpix({addrpix_0[388],addrpix_0[132]}));
	pe #(.ADR_WIDTH(2)) pe_0_133 (.state(state_0[535:532]),.ctrlreset(ctrlreset_0[535:532]),.reset(reset_0[535:532]),.enable(enable_0[133]),.valid(valid_0[133]),.rdpix(rdpix_0[133]),.addrpix({addrpix_0[389],addrpix_0[133]}));
	pe #(.ADR_WIDTH(2)) pe_0_134 (.state(state_0[539:536]),.ctrlreset(ctrlreset_0[539:536]),.reset(reset_0[539:536]),.enable(enable_0[134]),.valid(valid_0[134]),.rdpix(rdpix_0[134]),.addrpix({addrpix_0[390],addrpix_0[134]}));
	pe #(.ADR_WIDTH(2)) pe_0_135 (.state(state_0[543:540]),.ctrlreset(ctrlreset_0[543:540]),.reset(reset_0[543:540]),.enable(enable_0[135]),.valid(valid_0[135]),.rdpix(rdpix_0[135]),.addrpix({addrpix_0[391],addrpix_0[135]}));
	pe #(.ADR_WIDTH(2)) pe_0_136 (.state(state_0[547:544]),.ctrlreset(ctrlreset_0[547:544]),.reset(reset_0[547:544]),.enable(enable_0[136]),.valid(valid_0[136]),.rdpix(rdpix_0[136]),.addrpix({addrpix_0[392],addrpix_0[136]}));
	pe #(.ADR_WIDTH(2)) pe_0_137 (.state(state_0[551:548]),.ctrlreset(ctrlreset_0[551:548]),.reset(reset_0[551:548]),.enable(enable_0[137]),.valid(valid_0[137]),.rdpix(rdpix_0[137]),.addrpix({addrpix_0[393],addrpix_0[137]}));
	pe #(.ADR_WIDTH(2)) pe_0_138 (.state(state_0[555:552]),.ctrlreset(ctrlreset_0[555:552]),.reset(reset_0[555:552]),.enable(enable_0[138]),.valid(valid_0[138]),.rdpix(rdpix_0[138]),.addrpix({addrpix_0[394],addrpix_0[138]}));
	pe #(.ADR_WIDTH(2)) pe_0_139 (.state(state_0[559:556]),.ctrlreset(ctrlreset_0[559:556]),.reset(reset_0[559:556]),.enable(enable_0[139]),.valid(valid_0[139]),.rdpix(rdpix_0[139]),.addrpix({addrpix_0[395],addrpix_0[139]}));
	pe #(.ADR_WIDTH(2)) pe_0_140 (.state(state_0[563:560]),.ctrlreset(ctrlreset_0[563:560]),.reset(reset_0[563:560]),.enable(enable_0[140]),.valid(valid_0[140]),.rdpix(rdpix_0[140]),.addrpix({addrpix_0[396],addrpix_0[140]}));
	pe #(.ADR_WIDTH(2)) pe_0_141 (.state(state_0[567:564]),.ctrlreset(ctrlreset_0[567:564]),.reset(reset_0[567:564]),.enable(enable_0[141]),.valid(valid_0[141]),.rdpix(rdpix_0[141]),.addrpix({addrpix_0[397],addrpix_0[141]}));
	pe #(.ADR_WIDTH(2)) pe_0_142 (.state(state_0[571:568]),.ctrlreset(ctrlreset_0[571:568]),.reset(reset_0[571:568]),.enable(enable_0[142]),.valid(valid_0[142]),.rdpix(rdpix_0[142]),.addrpix({addrpix_0[398],addrpix_0[142]}));
	pe #(.ADR_WIDTH(2)) pe_0_143 (.state(state_0[575:572]),.ctrlreset(ctrlreset_0[575:572]),.reset(reset_0[575:572]),.enable(enable_0[143]),.valid(valid_0[143]),.rdpix(rdpix_0[143]),.addrpix({addrpix_0[399],addrpix_0[143]}));
	pe #(.ADR_WIDTH(2)) pe_0_144 (.state(state_0[579:576]),.ctrlreset(ctrlreset_0[579:576]),.reset(reset_0[579:576]),.enable(enable_0[144]),.valid(valid_0[144]),.rdpix(rdpix_0[144]),.addrpix({addrpix_0[400],addrpix_0[144]}));
	pe #(.ADR_WIDTH(2)) pe_0_145 (.state(state_0[583:580]),.ctrlreset(ctrlreset_0[583:580]),.reset(reset_0[583:580]),.enable(enable_0[145]),.valid(valid_0[145]),.rdpix(rdpix_0[145]),.addrpix({addrpix_0[401],addrpix_0[145]}));
	pe #(.ADR_WIDTH(2)) pe_0_146 (.state(state_0[587:584]),.ctrlreset(ctrlreset_0[587:584]),.reset(reset_0[587:584]),.enable(enable_0[146]),.valid(valid_0[146]),.rdpix(rdpix_0[146]),.addrpix({addrpix_0[402],addrpix_0[146]}));
	pe #(.ADR_WIDTH(2)) pe_0_147 (.state(state_0[591:588]),.ctrlreset(ctrlreset_0[591:588]),.reset(reset_0[591:588]),.enable(enable_0[147]),.valid(valid_0[147]),.rdpix(rdpix_0[147]),.addrpix({addrpix_0[403],addrpix_0[147]}));
	pe #(.ADR_WIDTH(2)) pe_0_148 (.state(state_0[595:592]),.ctrlreset(ctrlreset_0[595:592]),.reset(reset_0[595:592]),.enable(enable_0[148]),.valid(valid_0[148]),.rdpix(rdpix_0[148]),.addrpix({addrpix_0[404],addrpix_0[148]}));
	pe #(.ADR_WIDTH(2)) pe_0_149 (.state(state_0[599:596]),.ctrlreset(ctrlreset_0[599:596]),.reset(reset_0[599:596]),.enable(enable_0[149]),.valid(valid_0[149]),.rdpix(rdpix_0[149]),.addrpix({addrpix_0[405],addrpix_0[149]}));
	pe #(.ADR_WIDTH(2)) pe_0_150 (.state(state_0[603:600]),.ctrlreset(ctrlreset_0[603:600]),.reset(reset_0[603:600]),.enable(enable_0[150]),.valid(valid_0[150]),.rdpix(rdpix_0[150]),.addrpix({addrpix_0[406],addrpix_0[150]}));
	pe #(.ADR_WIDTH(2)) pe_0_151 (.state(state_0[607:604]),.ctrlreset(ctrlreset_0[607:604]),.reset(reset_0[607:604]),.enable(enable_0[151]),.valid(valid_0[151]),.rdpix(rdpix_0[151]),.addrpix({addrpix_0[407],addrpix_0[151]}));
	pe #(.ADR_WIDTH(2)) pe_0_152 (.state(state_0[611:608]),.ctrlreset(ctrlreset_0[611:608]),.reset(reset_0[611:608]),.enable(enable_0[152]),.valid(valid_0[152]),.rdpix(rdpix_0[152]),.addrpix({addrpix_0[408],addrpix_0[152]}));
	pe #(.ADR_WIDTH(2)) pe_0_153 (.state(state_0[615:612]),.ctrlreset(ctrlreset_0[615:612]),.reset(reset_0[615:612]),.enable(enable_0[153]),.valid(valid_0[153]),.rdpix(rdpix_0[153]),.addrpix({addrpix_0[409],addrpix_0[153]}));
	pe #(.ADR_WIDTH(2)) pe_0_154 (.state(state_0[619:616]),.ctrlreset(ctrlreset_0[619:616]),.reset(reset_0[619:616]),.enable(enable_0[154]),.valid(valid_0[154]),.rdpix(rdpix_0[154]),.addrpix({addrpix_0[410],addrpix_0[154]}));
	pe #(.ADR_WIDTH(2)) pe_0_155 (.state(state_0[623:620]),.ctrlreset(ctrlreset_0[623:620]),.reset(reset_0[623:620]),.enable(enable_0[155]),.valid(valid_0[155]),.rdpix(rdpix_0[155]),.addrpix({addrpix_0[411],addrpix_0[155]}));
	pe #(.ADR_WIDTH(2)) pe_0_156 (.state(state_0[627:624]),.ctrlreset(ctrlreset_0[627:624]),.reset(reset_0[627:624]),.enable(enable_0[156]),.valid(valid_0[156]),.rdpix(rdpix_0[156]),.addrpix({addrpix_0[412],addrpix_0[156]}));
	pe #(.ADR_WIDTH(2)) pe_0_157 (.state(state_0[631:628]),.ctrlreset(ctrlreset_0[631:628]),.reset(reset_0[631:628]),.enable(enable_0[157]),.valid(valid_0[157]),.rdpix(rdpix_0[157]),.addrpix({addrpix_0[413],addrpix_0[157]}));
	pe #(.ADR_WIDTH(2)) pe_0_158 (.state(state_0[635:632]),.ctrlreset(ctrlreset_0[635:632]),.reset(reset_0[635:632]),.enable(enable_0[158]),.valid(valid_0[158]),.rdpix(rdpix_0[158]),.addrpix({addrpix_0[414],addrpix_0[158]}));
	pe #(.ADR_WIDTH(2)) pe_0_159 (.state(state_0[639:636]),.ctrlreset(ctrlreset_0[639:636]),.reset(reset_0[639:636]),.enable(enable_0[159]),.valid(valid_0[159]),.rdpix(rdpix_0[159]),.addrpix({addrpix_0[415],addrpix_0[159]}));
	pe #(.ADR_WIDTH(2)) pe_0_160 (.state(state_0[643:640]),.ctrlreset(ctrlreset_0[643:640]),.reset(reset_0[643:640]),.enable(enable_0[160]),.valid(valid_0[160]),.rdpix(rdpix_0[160]),.addrpix({addrpix_0[416],addrpix_0[160]}));
	pe #(.ADR_WIDTH(2)) pe_0_161 (.state(state_0[647:644]),.ctrlreset(ctrlreset_0[647:644]),.reset(reset_0[647:644]),.enable(enable_0[161]),.valid(valid_0[161]),.rdpix(rdpix_0[161]),.addrpix({addrpix_0[417],addrpix_0[161]}));
	pe #(.ADR_WIDTH(2)) pe_0_162 (.state(state_0[651:648]),.ctrlreset(ctrlreset_0[651:648]),.reset(reset_0[651:648]),.enable(enable_0[162]),.valid(valid_0[162]),.rdpix(rdpix_0[162]),.addrpix({addrpix_0[418],addrpix_0[162]}));
	pe #(.ADR_WIDTH(2)) pe_0_163 (.state(state_0[655:652]),.ctrlreset(ctrlreset_0[655:652]),.reset(reset_0[655:652]),.enable(enable_0[163]),.valid(valid_0[163]),.rdpix(rdpix_0[163]),.addrpix({addrpix_0[419],addrpix_0[163]}));
	pe #(.ADR_WIDTH(2)) pe_0_164 (.state(state_0[659:656]),.ctrlreset(ctrlreset_0[659:656]),.reset(reset_0[659:656]),.enable(enable_0[164]),.valid(valid_0[164]),.rdpix(rdpix_0[164]),.addrpix({addrpix_0[420],addrpix_0[164]}));
	pe #(.ADR_WIDTH(2)) pe_0_165 (.state(state_0[663:660]),.ctrlreset(ctrlreset_0[663:660]),.reset(reset_0[663:660]),.enable(enable_0[165]),.valid(valid_0[165]),.rdpix(rdpix_0[165]),.addrpix({addrpix_0[421],addrpix_0[165]}));
	pe #(.ADR_WIDTH(2)) pe_0_166 (.state(state_0[667:664]),.ctrlreset(ctrlreset_0[667:664]),.reset(reset_0[667:664]),.enable(enable_0[166]),.valid(valid_0[166]),.rdpix(rdpix_0[166]),.addrpix({addrpix_0[422],addrpix_0[166]}));
	pe #(.ADR_WIDTH(2)) pe_0_167 (.state(state_0[671:668]),.ctrlreset(ctrlreset_0[671:668]),.reset(reset_0[671:668]),.enable(enable_0[167]),.valid(valid_0[167]),.rdpix(rdpix_0[167]),.addrpix({addrpix_0[423],addrpix_0[167]}));
	pe #(.ADR_WIDTH(2)) pe_0_168 (.state(state_0[675:672]),.ctrlreset(ctrlreset_0[675:672]),.reset(reset_0[675:672]),.enable(enable_0[168]),.valid(valid_0[168]),.rdpix(rdpix_0[168]),.addrpix({addrpix_0[424],addrpix_0[168]}));
	pe #(.ADR_WIDTH(2)) pe_0_169 (.state(state_0[679:676]),.ctrlreset(ctrlreset_0[679:676]),.reset(reset_0[679:676]),.enable(enable_0[169]),.valid(valid_0[169]),.rdpix(rdpix_0[169]),.addrpix({addrpix_0[425],addrpix_0[169]}));
	pe #(.ADR_WIDTH(2)) pe_0_170 (.state(state_0[683:680]),.ctrlreset(ctrlreset_0[683:680]),.reset(reset_0[683:680]),.enable(enable_0[170]),.valid(valid_0[170]),.rdpix(rdpix_0[170]),.addrpix({addrpix_0[426],addrpix_0[170]}));
	pe #(.ADR_WIDTH(2)) pe_0_171 (.state(state_0[687:684]),.ctrlreset(ctrlreset_0[687:684]),.reset(reset_0[687:684]),.enable(enable_0[171]),.valid(valid_0[171]),.rdpix(rdpix_0[171]),.addrpix({addrpix_0[427],addrpix_0[171]}));
	pe #(.ADR_WIDTH(2)) pe_0_172 (.state(state_0[691:688]),.ctrlreset(ctrlreset_0[691:688]),.reset(reset_0[691:688]),.enable(enable_0[172]),.valid(valid_0[172]),.rdpix(rdpix_0[172]),.addrpix({addrpix_0[428],addrpix_0[172]}));
	pe #(.ADR_WIDTH(2)) pe_0_173 (.state(state_0[695:692]),.ctrlreset(ctrlreset_0[695:692]),.reset(reset_0[695:692]),.enable(enable_0[173]),.valid(valid_0[173]),.rdpix(rdpix_0[173]),.addrpix({addrpix_0[429],addrpix_0[173]}));
	pe #(.ADR_WIDTH(2)) pe_0_174 (.state(state_0[699:696]),.ctrlreset(ctrlreset_0[699:696]),.reset(reset_0[699:696]),.enable(enable_0[174]),.valid(valid_0[174]),.rdpix(rdpix_0[174]),.addrpix({addrpix_0[430],addrpix_0[174]}));
	pe #(.ADR_WIDTH(2)) pe_0_175 (.state(state_0[703:700]),.ctrlreset(ctrlreset_0[703:700]),.reset(reset_0[703:700]),.enable(enable_0[175]),.valid(valid_0[175]),.rdpix(rdpix_0[175]),.addrpix({addrpix_0[431],addrpix_0[175]}));
	pe #(.ADR_WIDTH(2)) pe_0_176 (.state(state_0[707:704]),.ctrlreset(ctrlreset_0[707:704]),.reset(reset_0[707:704]),.enable(enable_0[176]),.valid(valid_0[176]),.rdpix(rdpix_0[176]),.addrpix({addrpix_0[432],addrpix_0[176]}));
	pe #(.ADR_WIDTH(2)) pe_0_177 (.state(state_0[711:708]),.ctrlreset(ctrlreset_0[711:708]),.reset(reset_0[711:708]),.enable(enable_0[177]),.valid(valid_0[177]),.rdpix(rdpix_0[177]),.addrpix({addrpix_0[433],addrpix_0[177]}));
	pe #(.ADR_WIDTH(2)) pe_0_178 (.state(state_0[715:712]),.ctrlreset(ctrlreset_0[715:712]),.reset(reset_0[715:712]),.enable(enable_0[178]),.valid(valid_0[178]),.rdpix(rdpix_0[178]),.addrpix({addrpix_0[434],addrpix_0[178]}));
	pe #(.ADR_WIDTH(2)) pe_0_179 (.state(state_0[719:716]),.ctrlreset(ctrlreset_0[719:716]),.reset(reset_0[719:716]),.enable(enable_0[179]),.valid(valid_0[179]),.rdpix(rdpix_0[179]),.addrpix({addrpix_0[435],addrpix_0[179]}));
	pe #(.ADR_WIDTH(2)) pe_0_180 (.state(state_0[723:720]),.ctrlreset(ctrlreset_0[723:720]),.reset(reset_0[723:720]),.enable(enable_0[180]),.valid(valid_0[180]),.rdpix(rdpix_0[180]),.addrpix({addrpix_0[436],addrpix_0[180]}));
	pe #(.ADR_WIDTH(2)) pe_0_181 (.state(state_0[727:724]),.ctrlreset(ctrlreset_0[727:724]),.reset(reset_0[727:724]),.enable(enable_0[181]),.valid(valid_0[181]),.rdpix(rdpix_0[181]),.addrpix({addrpix_0[437],addrpix_0[181]}));
	pe #(.ADR_WIDTH(2)) pe_0_182 (.state(state_0[731:728]),.ctrlreset(ctrlreset_0[731:728]),.reset(reset_0[731:728]),.enable(enable_0[182]),.valid(valid_0[182]),.rdpix(rdpix_0[182]),.addrpix({addrpix_0[438],addrpix_0[182]}));
	pe #(.ADR_WIDTH(2)) pe_0_183 (.state(state_0[735:732]),.ctrlreset(ctrlreset_0[735:732]),.reset(reset_0[735:732]),.enable(enable_0[183]),.valid(valid_0[183]),.rdpix(rdpix_0[183]),.addrpix({addrpix_0[439],addrpix_0[183]}));
	pe #(.ADR_WIDTH(2)) pe_0_184 (.state(state_0[739:736]),.ctrlreset(ctrlreset_0[739:736]),.reset(reset_0[739:736]),.enable(enable_0[184]),.valid(valid_0[184]),.rdpix(rdpix_0[184]),.addrpix({addrpix_0[440],addrpix_0[184]}));
	pe #(.ADR_WIDTH(2)) pe_0_185 (.state(state_0[743:740]),.ctrlreset(ctrlreset_0[743:740]),.reset(reset_0[743:740]),.enable(enable_0[185]),.valid(valid_0[185]),.rdpix(rdpix_0[185]),.addrpix({addrpix_0[441],addrpix_0[185]}));
	pe #(.ADR_WIDTH(2)) pe_0_186 (.state(state_0[747:744]),.ctrlreset(ctrlreset_0[747:744]),.reset(reset_0[747:744]),.enable(enable_0[186]),.valid(valid_0[186]),.rdpix(rdpix_0[186]),.addrpix({addrpix_0[442],addrpix_0[186]}));
	pe #(.ADR_WIDTH(2)) pe_0_187 (.state(state_0[751:748]),.ctrlreset(ctrlreset_0[751:748]),.reset(reset_0[751:748]),.enable(enable_0[187]),.valid(valid_0[187]),.rdpix(rdpix_0[187]),.addrpix({addrpix_0[443],addrpix_0[187]}));
	pe #(.ADR_WIDTH(2)) pe_0_188 (.state(state_0[755:752]),.ctrlreset(ctrlreset_0[755:752]),.reset(reset_0[755:752]),.enable(enable_0[188]),.valid(valid_0[188]),.rdpix(rdpix_0[188]),.addrpix({addrpix_0[444],addrpix_0[188]}));
	pe #(.ADR_WIDTH(2)) pe_0_189 (.state(state_0[759:756]),.ctrlreset(ctrlreset_0[759:756]),.reset(reset_0[759:756]),.enable(enable_0[189]),.valid(valid_0[189]),.rdpix(rdpix_0[189]),.addrpix({addrpix_0[445],addrpix_0[189]}));
	pe #(.ADR_WIDTH(2)) pe_0_190 (.state(state_0[763:760]),.ctrlreset(ctrlreset_0[763:760]),.reset(reset_0[763:760]),.enable(enable_0[190]),.valid(valid_0[190]),.rdpix(rdpix_0[190]),.addrpix({addrpix_0[446],addrpix_0[190]}));
	pe #(.ADR_WIDTH(2)) pe_0_191 (.state(state_0[767:764]),.ctrlreset(ctrlreset_0[767:764]),.reset(reset_0[767:764]),.enable(enable_0[191]),.valid(valid_0[191]),.rdpix(rdpix_0[191]),.addrpix({addrpix_0[447],addrpix_0[191]}));
	pe #(.ADR_WIDTH(2)) pe_0_192 (.state(state_0[771:768]),.ctrlreset(ctrlreset_0[771:768]),.reset(reset_0[771:768]),.enable(enable_0[192]),.valid(valid_0[192]),.rdpix(rdpix_0[192]),.addrpix({addrpix_0[448],addrpix_0[192]}));
	pe #(.ADR_WIDTH(2)) pe_0_193 (.state(state_0[775:772]),.ctrlreset(ctrlreset_0[775:772]),.reset(reset_0[775:772]),.enable(enable_0[193]),.valid(valid_0[193]),.rdpix(rdpix_0[193]),.addrpix({addrpix_0[449],addrpix_0[193]}));
	pe #(.ADR_WIDTH(2)) pe_0_194 (.state(state_0[779:776]),.ctrlreset(ctrlreset_0[779:776]),.reset(reset_0[779:776]),.enable(enable_0[194]),.valid(valid_0[194]),.rdpix(rdpix_0[194]),.addrpix({addrpix_0[450],addrpix_0[194]}));
	pe #(.ADR_WIDTH(2)) pe_0_195 (.state(state_0[783:780]),.ctrlreset(ctrlreset_0[783:780]),.reset(reset_0[783:780]),.enable(enable_0[195]),.valid(valid_0[195]),.rdpix(rdpix_0[195]),.addrpix({addrpix_0[451],addrpix_0[195]}));
	pe #(.ADR_WIDTH(2)) pe_0_196 (.state(state_0[787:784]),.ctrlreset(ctrlreset_0[787:784]),.reset(reset_0[787:784]),.enable(enable_0[196]),.valid(valid_0[196]),.rdpix(rdpix_0[196]),.addrpix({addrpix_0[452],addrpix_0[196]}));
	pe #(.ADR_WIDTH(2)) pe_0_197 (.state(state_0[791:788]),.ctrlreset(ctrlreset_0[791:788]),.reset(reset_0[791:788]),.enable(enable_0[197]),.valid(valid_0[197]),.rdpix(rdpix_0[197]),.addrpix({addrpix_0[453],addrpix_0[197]}));
	pe #(.ADR_WIDTH(2)) pe_0_198 (.state(state_0[795:792]),.ctrlreset(ctrlreset_0[795:792]),.reset(reset_0[795:792]),.enable(enable_0[198]),.valid(valid_0[198]),.rdpix(rdpix_0[198]),.addrpix({addrpix_0[454],addrpix_0[198]}));
	pe #(.ADR_WIDTH(2)) pe_0_199 (.state(state_0[799:796]),.ctrlreset(ctrlreset_0[799:796]),.reset(reset_0[799:796]),.enable(enable_0[199]),.valid(valid_0[199]),.rdpix(rdpix_0[199]),.addrpix({addrpix_0[455],addrpix_0[199]}));
	pe #(.ADR_WIDTH(2)) pe_0_200 (.state(state_0[803:800]),.ctrlreset(ctrlreset_0[803:800]),.reset(reset_0[803:800]),.enable(enable_0[200]),.valid(valid_0[200]),.rdpix(rdpix_0[200]),.addrpix({addrpix_0[456],addrpix_0[200]}));
	pe #(.ADR_WIDTH(2)) pe_0_201 (.state(state_0[807:804]),.ctrlreset(ctrlreset_0[807:804]),.reset(reset_0[807:804]),.enable(enable_0[201]),.valid(valid_0[201]),.rdpix(rdpix_0[201]),.addrpix({addrpix_0[457],addrpix_0[201]}));
	pe #(.ADR_WIDTH(2)) pe_0_202 (.state(state_0[811:808]),.ctrlreset(ctrlreset_0[811:808]),.reset(reset_0[811:808]),.enable(enable_0[202]),.valid(valid_0[202]),.rdpix(rdpix_0[202]),.addrpix({addrpix_0[458],addrpix_0[202]}));
	pe #(.ADR_WIDTH(2)) pe_0_203 (.state(state_0[815:812]),.ctrlreset(ctrlreset_0[815:812]),.reset(reset_0[815:812]),.enable(enable_0[203]),.valid(valid_0[203]),.rdpix(rdpix_0[203]),.addrpix({addrpix_0[459],addrpix_0[203]}));
	pe #(.ADR_WIDTH(2)) pe_0_204 (.state(state_0[819:816]),.ctrlreset(ctrlreset_0[819:816]),.reset(reset_0[819:816]),.enable(enable_0[204]),.valid(valid_0[204]),.rdpix(rdpix_0[204]),.addrpix({addrpix_0[460],addrpix_0[204]}));
	pe #(.ADR_WIDTH(2)) pe_0_205 (.state(state_0[823:820]),.ctrlreset(ctrlreset_0[823:820]),.reset(reset_0[823:820]),.enable(enable_0[205]),.valid(valid_0[205]),.rdpix(rdpix_0[205]),.addrpix({addrpix_0[461],addrpix_0[205]}));
	pe #(.ADR_WIDTH(2)) pe_0_206 (.state(state_0[827:824]),.ctrlreset(ctrlreset_0[827:824]),.reset(reset_0[827:824]),.enable(enable_0[206]),.valid(valid_0[206]),.rdpix(rdpix_0[206]),.addrpix({addrpix_0[462],addrpix_0[206]}));
	pe #(.ADR_WIDTH(2)) pe_0_207 (.state(state_0[831:828]),.ctrlreset(ctrlreset_0[831:828]),.reset(reset_0[831:828]),.enable(enable_0[207]),.valid(valid_0[207]),.rdpix(rdpix_0[207]),.addrpix({addrpix_0[463],addrpix_0[207]}));
	pe #(.ADR_WIDTH(2)) pe_0_208 (.state(state_0[835:832]),.ctrlreset(ctrlreset_0[835:832]),.reset(reset_0[835:832]),.enable(enable_0[208]),.valid(valid_0[208]),.rdpix(rdpix_0[208]),.addrpix({addrpix_0[464],addrpix_0[208]}));
	pe #(.ADR_WIDTH(2)) pe_0_209 (.state(state_0[839:836]),.ctrlreset(ctrlreset_0[839:836]),.reset(reset_0[839:836]),.enable(enable_0[209]),.valid(valid_0[209]),.rdpix(rdpix_0[209]),.addrpix({addrpix_0[465],addrpix_0[209]}));
	pe #(.ADR_WIDTH(2)) pe_0_210 (.state(state_0[843:840]),.ctrlreset(ctrlreset_0[843:840]),.reset(reset_0[843:840]),.enable(enable_0[210]),.valid(valid_0[210]),.rdpix(rdpix_0[210]),.addrpix({addrpix_0[466],addrpix_0[210]}));
	pe #(.ADR_WIDTH(2)) pe_0_211 (.state(state_0[847:844]),.ctrlreset(ctrlreset_0[847:844]),.reset(reset_0[847:844]),.enable(enable_0[211]),.valid(valid_0[211]),.rdpix(rdpix_0[211]),.addrpix({addrpix_0[467],addrpix_0[211]}));
	pe #(.ADR_WIDTH(2)) pe_0_212 (.state(state_0[851:848]),.ctrlreset(ctrlreset_0[851:848]),.reset(reset_0[851:848]),.enable(enable_0[212]),.valid(valid_0[212]),.rdpix(rdpix_0[212]),.addrpix({addrpix_0[468],addrpix_0[212]}));
	pe #(.ADR_WIDTH(2)) pe_0_213 (.state(state_0[855:852]),.ctrlreset(ctrlreset_0[855:852]),.reset(reset_0[855:852]),.enable(enable_0[213]),.valid(valid_0[213]),.rdpix(rdpix_0[213]),.addrpix({addrpix_0[469],addrpix_0[213]}));
	pe #(.ADR_WIDTH(2)) pe_0_214 (.state(state_0[859:856]),.ctrlreset(ctrlreset_0[859:856]),.reset(reset_0[859:856]),.enable(enable_0[214]),.valid(valid_0[214]),.rdpix(rdpix_0[214]),.addrpix({addrpix_0[470],addrpix_0[214]}));
	pe #(.ADR_WIDTH(2)) pe_0_215 (.state(state_0[863:860]),.ctrlreset(ctrlreset_0[863:860]),.reset(reset_0[863:860]),.enable(enable_0[215]),.valid(valid_0[215]),.rdpix(rdpix_0[215]),.addrpix({addrpix_0[471],addrpix_0[215]}));
	pe #(.ADR_WIDTH(2)) pe_0_216 (.state(state_0[867:864]),.ctrlreset(ctrlreset_0[867:864]),.reset(reset_0[867:864]),.enable(enable_0[216]),.valid(valid_0[216]),.rdpix(rdpix_0[216]),.addrpix({addrpix_0[472],addrpix_0[216]}));
	pe #(.ADR_WIDTH(2)) pe_0_217 (.state(state_0[871:868]),.ctrlreset(ctrlreset_0[871:868]),.reset(reset_0[871:868]),.enable(enable_0[217]),.valid(valid_0[217]),.rdpix(rdpix_0[217]),.addrpix({addrpix_0[473],addrpix_0[217]}));
	pe #(.ADR_WIDTH(2)) pe_0_218 (.state(state_0[875:872]),.ctrlreset(ctrlreset_0[875:872]),.reset(reset_0[875:872]),.enable(enable_0[218]),.valid(valid_0[218]),.rdpix(rdpix_0[218]),.addrpix({addrpix_0[474],addrpix_0[218]}));
	pe #(.ADR_WIDTH(2)) pe_0_219 (.state(state_0[879:876]),.ctrlreset(ctrlreset_0[879:876]),.reset(reset_0[879:876]),.enable(enable_0[219]),.valid(valid_0[219]),.rdpix(rdpix_0[219]),.addrpix({addrpix_0[475],addrpix_0[219]}));
	pe #(.ADR_WIDTH(2)) pe_0_220 (.state(state_0[883:880]),.ctrlreset(ctrlreset_0[883:880]),.reset(reset_0[883:880]),.enable(enable_0[220]),.valid(valid_0[220]),.rdpix(rdpix_0[220]),.addrpix({addrpix_0[476],addrpix_0[220]}));
	pe #(.ADR_WIDTH(2)) pe_0_221 (.state(state_0[887:884]),.ctrlreset(ctrlreset_0[887:884]),.reset(reset_0[887:884]),.enable(enable_0[221]),.valid(valid_0[221]),.rdpix(rdpix_0[221]),.addrpix({addrpix_0[477],addrpix_0[221]}));
	pe #(.ADR_WIDTH(2)) pe_0_222 (.state(state_0[891:888]),.ctrlreset(ctrlreset_0[891:888]),.reset(reset_0[891:888]),.enable(enable_0[222]),.valid(valid_0[222]),.rdpix(rdpix_0[222]),.addrpix({addrpix_0[478],addrpix_0[222]}));
	pe #(.ADR_WIDTH(2)) pe_0_223 (.state(state_0[895:892]),.ctrlreset(ctrlreset_0[895:892]),.reset(reset_0[895:892]),.enable(enable_0[223]),.valid(valid_0[223]),.rdpix(rdpix_0[223]),.addrpix({addrpix_0[479],addrpix_0[223]}));
	pe #(.ADR_WIDTH(2)) pe_0_224 (.state(state_0[899:896]),.ctrlreset(ctrlreset_0[899:896]),.reset(reset_0[899:896]),.enable(enable_0[224]),.valid(valid_0[224]),.rdpix(rdpix_0[224]),.addrpix({addrpix_0[480],addrpix_0[224]}));
	pe #(.ADR_WIDTH(2)) pe_0_225 (.state(state_0[903:900]),.ctrlreset(ctrlreset_0[903:900]),.reset(reset_0[903:900]),.enable(enable_0[225]),.valid(valid_0[225]),.rdpix(rdpix_0[225]),.addrpix({addrpix_0[481],addrpix_0[225]}));
	pe #(.ADR_WIDTH(2)) pe_0_226 (.state(state_0[907:904]),.ctrlreset(ctrlreset_0[907:904]),.reset(reset_0[907:904]),.enable(enable_0[226]),.valid(valid_0[226]),.rdpix(rdpix_0[226]),.addrpix({addrpix_0[482],addrpix_0[226]}));
	pe #(.ADR_WIDTH(2)) pe_0_227 (.state(state_0[911:908]),.ctrlreset(ctrlreset_0[911:908]),.reset(reset_0[911:908]),.enable(enable_0[227]),.valid(valid_0[227]),.rdpix(rdpix_0[227]),.addrpix({addrpix_0[483],addrpix_0[227]}));
	pe #(.ADR_WIDTH(2)) pe_0_228 (.state(state_0[915:912]),.ctrlreset(ctrlreset_0[915:912]),.reset(reset_0[915:912]),.enable(enable_0[228]),.valid(valid_0[228]),.rdpix(rdpix_0[228]),.addrpix({addrpix_0[484],addrpix_0[228]}));
	pe #(.ADR_WIDTH(2)) pe_0_229 (.state(state_0[919:916]),.ctrlreset(ctrlreset_0[919:916]),.reset(reset_0[919:916]),.enable(enable_0[229]),.valid(valid_0[229]),.rdpix(rdpix_0[229]),.addrpix({addrpix_0[485],addrpix_0[229]}));
	pe #(.ADR_WIDTH(2)) pe_0_230 (.state(state_0[923:920]),.ctrlreset(ctrlreset_0[923:920]),.reset(reset_0[923:920]),.enable(enable_0[230]),.valid(valid_0[230]),.rdpix(rdpix_0[230]),.addrpix({addrpix_0[486],addrpix_0[230]}));
	pe #(.ADR_WIDTH(2)) pe_0_231 (.state(state_0[927:924]),.ctrlreset(ctrlreset_0[927:924]),.reset(reset_0[927:924]),.enable(enable_0[231]),.valid(valid_0[231]),.rdpix(rdpix_0[231]),.addrpix({addrpix_0[487],addrpix_0[231]}));
	pe #(.ADR_WIDTH(2)) pe_0_232 (.state(state_0[931:928]),.ctrlreset(ctrlreset_0[931:928]),.reset(reset_0[931:928]),.enable(enable_0[232]),.valid(valid_0[232]),.rdpix(rdpix_0[232]),.addrpix({addrpix_0[488],addrpix_0[232]}));
	pe #(.ADR_WIDTH(2)) pe_0_233 (.state(state_0[935:932]),.ctrlreset(ctrlreset_0[935:932]),.reset(reset_0[935:932]),.enable(enable_0[233]),.valid(valid_0[233]),.rdpix(rdpix_0[233]),.addrpix({addrpix_0[489],addrpix_0[233]}));
	pe #(.ADR_WIDTH(2)) pe_0_234 (.state(state_0[939:936]),.ctrlreset(ctrlreset_0[939:936]),.reset(reset_0[939:936]),.enable(enable_0[234]),.valid(valid_0[234]),.rdpix(rdpix_0[234]),.addrpix({addrpix_0[490],addrpix_0[234]}));
	pe #(.ADR_WIDTH(2)) pe_0_235 (.state(state_0[943:940]),.ctrlreset(ctrlreset_0[943:940]),.reset(reset_0[943:940]),.enable(enable_0[235]),.valid(valid_0[235]),.rdpix(rdpix_0[235]),.addrpix({addrpix_0[491],addrpix_0[235]}));
	pe #(.ADR_WIDTH(2)) pe_0_236 (.state(state_0[947:944]),.ctrlreset(ctrlreset_0[947:944]),.reset(reset_0[947:944]),.enable(enable_0[236]),.valid(valid_0[236]),.rdpix(rdpix_0[236]),.addrpix({addrpix_0[492],addrpix_0[236]}));
	pe #(.ADR_WIDTH(2)) pe_0_237 (.state(state_0[951:948]),.ctrlreset(ctrlreset_0[951:948]),.reset(reset_0[951:948]),.enable(enable_0[237]),.valid(valid_0[237]),.rdpix(rdpix_0[237]),.addrpix({addrpix_0[493],addrpix_0[237]}));
	pe #(.ADR_WIDTH(2)) pe_0_238 (.state(state_0[955:952]),.ctrlreset(ctrlreset_0[955:952]),.reset(reset_0[955:952]),.enable(enable_0[238]),.valid(valid_0[238]),.rdpix(rdpix_0[238]),.addrpix({addrpix_0[494],addrpix_0[238]}));
	pe #(.ADR_WIDTH(2)) pe_0_239 (.state(state_0[959:956]),.ctrlreset(ctrlreset_0[959:956]),.reset(reset_0[959:956]),.enable(enable_0[239]),.valid(valid_0[239]),.rdpix(rdpix_0[239]),.addrpix({addrpix_0[495],addrpix_0[239]}));
	pe #(.ADR_WIDTH(2)) pe_0_240 (.state(state_0[963:960]),.ctrlreset(ctrlreset_0[963:960]),.reset(reset_0[963:960]),.enable(enable_0[240]),.valid(valid_0[240]),.rdpix(rdpix_0[240]),.addrpix({addrpix_0[496],addrpix_0[240]}));
	pe #(.ADR_WIDTH(2)) pe_0_241 (.state(state_0[967:964]),.ctrlreset(ctrlreset_0[967:964]),.reset(reset_0[967:964]),.enable(enable_0[241]),.valid(valid_0[241]),.rdpix(rdpix_0[241]),.addrpix({addrpix_0[497],addrpix_0[241]}));
	pe #(.ADR_WIDTH(2)) pe_0_242 (.state(state_0[971:968]),.ctrlreset(ctrlreset_0[971:968]),.reset(reset_0[971:968]),.enable(enable_0[242]),.valid(valid_0[242]),.rdpix(rdpix_0[242]),.addrpix({addrpix_0[498],addrpix_0[242]}));
	pe #(.ADR_WIDTH(2)) pe_0_243 (.state(state_0[975:972]),.ctrlreset(ctrlreset_0[975:972]),.reset(reset_0[975:972]),.enable(enable_0[243]),.valid(valid_0[243]),.rdpix(rdpix_0[243]),.addrpix({addrpix_0[499],addrpix_0[243]}));
	pe #(.ADR_WIDTH(2)) pe_0_244 (.state(state_0[979:976]),.ctrlreset(ctrlreset_0[979:976]),.reset(reset_0[979:976]),.enable(enable_0[244]),.valid(valid_0[244]),.rdpix(rdpix_0[244]),.addrpix({addrpix_0[500],addrpix_0[244]}));
	pe #(.ADR_WIDTH(2)) pe_0_245 (.state(state_0[983:980]),.ctrlreset(ctrlreset_0[983:980]),.reset(reset_0[983:980]),.enable(enable_0[245]),.valid(valid_0[245]),.rdpix(rdpix_0[245]),.addrpix({addrpix_0[501],addrpix_0[245]}));
	pe #(.ADR_WIDTH(2)) pe_0_246 (.state(state_0[987:984]),.ctrlreset(ctrlreset_0[987:984]),.reset(reset_0[987:984]),.enable(enable_0[246]),.valid(valid_0[246]),.rdpix(rdpix_0[246]),.addrpix({addrpix_0[502],addrpix_0[246]}));
	pe #(.ADR_WIDTH(2)) pe_0_247 (.state(state_0[991:988]),.ctrlreset(ctrlreset_0[991:988]),.reset(reset_0[991:988]),.enable(enable_0[247]),.valid(valid_0[247]),.rdpix(rdpix_0[247]),.addrpix({addrpix_0[503],addrpix_0[247]}));
	pe #(.ADR_WIDTH(2)) pe_0_248 (.state(state_0[995:992]),.ctrlreset(ctrlreset_0[995:992]),.reset(reset_0[995:992]),.enable(enable_0[248]),.valid(valid_0[248]),.rdpix(rdpix_0[248]),.addrpix({addrpix_0[504],addrpix_0[248]}));
	pe #(.ADR_WIDTH(2)) pe_0_249 (.state(state_0[999:996]),.ctrlreset(ctrlreset_0[999:996]),.reset(reset_0[999:996]),.enable(enable_0[249]),.valid(valid_0[249]),.rdpix(rdpix_0[249]),.addrpix({addrpix_0[505],addrpix_0[249]}));
	pe #(.ADR_WIDTH(2)) pe_0_250 (.state(state_0[1003:1000]),.ctrlreset(ctrlreset_0[1003:1000]),.reset(reset_0[1003:1000]),.enable(enable_0[250]),.valid(valid_0[250]),.rdpix(rdpix_0[250]),.addrpix({addrpix_0[506],addrpix_0[250]}));
	pe #(.ADR_WIDTH(2)) pe_0_251 (.state(state_0[1007:1004]),.ctrlreset(ctrlreset_0[1007:1004]),.reset(reset_0[1007:1004]),.enable(enable_0[251]),.valid(valid_0[251]),.rdpix(rdpix_0[251]),.addrpix({addrpix_0[507],addrpix_0[251]}));
	pe #(.ADR_WIDTH(2)) pe_0_252 (.state(state_0[1011:1008]),.ctrlreset(ctrlreset_0[1011:1008]),.reset(reset_0[1011:1008]),.enable(enable_0[252]),.valid(valid_0[252]),.rdpix(rdpix_0[252]),.addrpix({addrpix_0[508],addrpix_0[252]}));
	pe #(.ADR_WIDTH(2)) pe_0_253 (.state(state_0[1015:1012]),.ctrlreset(ctrlreset_0[1015:1012]),.reset(reset_0[1015:1012]),.enable(enable_0[253]),.valid(valid_0[253]),.rdpix(rdpix_0[253]),.addrpix({addrpix_0[509],addrpix_0[253]}));
	pe #(.ADR_WIDTH(2)) pe_0_254 (.state(state_0[1019:1016]),.ctrlreset(ctrlreset_0[1019:1016]),.reset(reset_0[1019:1016]),.enable(enable_0[254]),.valid(valid_0[254]),.rdpix(rdpix_0[254]),.addrpix({addrpix_0[510],addrpix_0[254]}));
	pe #(.ADR_WIDTH(2)) pe_0_255 (.state(state_0[1023:1020]),.ctrlreset(ctrlreset_0[1023:1020]),.reset(reset_0[1023:1020]),.enable(enable_0[255]),.valid(valid_0[255]),.rdpix(rdpix_0[255]),.addrpix({addrpix_0[511],addrpix_0[255]}));
assign addrpix[1:0] = {|addrpix_0[511:256],|addrpix_0[255:0]};
// Level 1
wire [255:0] state_1;
wire [255:0] reset_1;
wire [255:0] ctrlreset_1;
wire [63:0] enable_1;
wire [63:0] rdpix_1;
wire [63:0] valid_1;
wire [127:0] addrpix_1;
	pe #(.ADR_WIDTH(2)) pe_1_0 (.state(state_1[3:0]),.ctrlreset(ctrlreset_1[3:0]),.reset(reset_1[3:0]),.enable(enable_1[0]),.valid(valid_1[0]),.rdpix(rdpix_1[0]),.addrpix({addrpix_1[64],addrpix_1[0]}));
	pe #(.ADR_WIDTH(2)) pe_1_1 (.state(state_1[7:4]),.ctrlreset(ctrlreset_1[7:4]),.reset(reset_1[7:4]),.enable(enable_1[1]),.valid(valid_1[1]),.rdpix(rdpix_1[1]),.addrpix({addrpix_1[65],addrpix_1[1]}));
	pe #(.ADR_WIDTH(2)) pe_1_2 (.state(state_1[11:8]),.ctrlreset(ctrlreset_1[11:8]),.reset(reset_1[11:8]),.enable(enable_1[2]),.valid(valid_1[2]),.rdpix(rdpix_1[2]),.addrpix({addrpix_1[66],addrpix_1[2]}));
	pe #(.ADR_WIDTH(2)) pe_1_3 (.state(state_1[15:12]),.ctrlreset(ctrlreset_1[15:12]),.reset(reset_1[15:12]),.enable(enable_1[3]),.valid(valid_1[3]),.rdpix(rdpix_1[3]),.addrpix({addrpix_1[67],addrpix_1[3]}));
	pe #(.ADR_WIDTH(2)) pe_1_4 (.state(state_1[19:16]),.ctrlreset(ctrlreset_1[19:16]),.reset(reset_1[19:16]),.enable(enable_1[4]),.valid(valid_1[4]),.rdpix(rdpix_1[4]),.addrpix({addrpix_1[68],addrpix_1[4]}));
	pe #(.ADR_WIDTH(2)) pe_1_5 (.state(state_1[23:20]),.ctrlreset(ctrlreset_1[23:20]),.reset(reset_1[23:20]),.enable(enable_1[5]),.valid(valid_1[5]),.rdpix(rdpix_1[5]),.addrpix({addrpix_1[69],addrpix_1[5]}));
	pe #(.ADR_WIDTH(2)) pe_1_6 (.state(state_1[27:24]),.ctrlreset(ctrlreset_1[27:24]),.reset(reset_1[27:24]),.enable(enable_1[6]),.valid(valid_1[6]),.rdpix(rdpix_1[6]),.addrpix({addrpix_1[70],addrpix_1[6]}));
	pe #(.ADR_WIDTH(2)) pe_1_7 (.state(state_1[31:28]),.ctrlreset(ctrlreset_1[31:28]),.reset(reset_1[31:28]),.enable(enable_1[7]),.valid(valid_1[7]),.rdpix(rdpix_1[7]),.addrpix({addrpix_1[71],addrpix_1[7]}));
	pe #(.ADR_WIDTH(2)) pe_1_8 (.state(state_1[35:32]),.ctrlreset(ctrlreset_1[35:32]),.reset(reset_1[35:32]),.enable(enable_1[8]),.valid(valid_1[8]),.rdpix(rdpix_1[8]),.addrpix({addrpix_1[72],addrpix_1[8]}));
	pe #(.ADR_WIDTH(2)) pe_1_9 (.state(state_1[39:36]),.ctrlreset(ctrlreset_1[39:36]),.reset(reset_1[39:36]),.enable(enable_1[9]),.valid(valid_1[9]),.rdpix(rdpix_1[9]),.addrpix({addrpix_1[73],addrpix_1[9]}));
	pe #(.ADR_WIDTH(2)) pe_1_10 (.state(state_1[43:40]),.ctrlreset(ctrlreset_1[43:40]),.reset(reset_1[43:40]),.enable(enable_1[10]),.valid(valid_1[10]),.rdpix(rdpix_1[10]),.addrpix({addrpix_1[74],addrpix_1[10]}));
	pe #(.ADR_WIDTH(2)) pe_1_11 (.state(state_1[47:44]),.ctrlreset(ctrlreset_1[47:44]),.reset(reset_1[47:44]),.enable(enable_1[11]),.valid(valid_1[11]),.rdpix(rdpix_1[11]),.addrpix({addrpix_1[75],addrpix_1[11]}));
	pe #(.ADR_WIDTH(2)) pe_1_12 (.state(state_1[51:48]),.ctrlreset(ctrlreset_1[51:48]),.reset(reset_1[51:48]),.enable(enable_1[12]),.valid(valid_1[12]),.rdpix(rdpix_1[12]),.addrpix({addrpix_1[76],addrpix_1[12]}));
	pe #(.ADR_WIDTH(2)) pe_1_13 (.state(state_1[55:52]),.ctrlreset(ctrlreset_1[55:52]),.reset(reset_1[55:52]),.enable(enable_1[13]),.valid(valid_1[13]),.rdpix(rdpix_1[13]),.addrpix({addrpix_1[77],addrpix_1[13]}));
	pe #(.ADR_WIDTH(2)) pe_1_14 (.state(state_1[59:56]),.ctrlreset(ctrlreset_1[59:56]),.reset(reset_1[59:56]),.enable(enable_1[14]),.valid(valid_1[14]),.rdpix(rdpix_1[14]),.addrpix({addrpix_1[78],addrpix_1[14]}));
	pe #(.ADR_WIDTH(2)) pe_1_15 (.state(state_1[63:60]),.ctrlreset(ctrlreset_1[63:60]),.reset(reset_1[63:60]),.enable(enable_1[15]),.valid(valid_1[15]),.rdpix(rdpix_1[15]),.addrpix({addrpix_1[79],addrpix_1[15]}));
	pe #(.ADR_WIDTH(2)) pe_1_16 (.state(state_1[67:64]),.ctrlreset(ctrlreset_1[67:64]),.reset(reset_1[67:64]),.enable(enable_1[16]),.valid(valid_1[16]),.rdpix(rdpix_1[16]),.addrpix({addrpix_1[80],addrpix_1[16]}));
	pe #(.ADR_WIDTH(2)) pe_1_17 (.state(state_1[71:68]),.ctrlreset(ctrlreset_1[71:68]),.reset(reset_1[71:68]),.enable(enable_1[17]),.valid(valid_1[17]),.rdpix(rdpix_1[17]),.addrpix({addrpix_1[81],addrpix_1[17]}));
	pe #(.ADR_WIDTH(2)) pe_1_18 (.state(state_1[75:72]),.ctrlreset(ctrlreset_1[75:72]),.reset(reset_1[75:72]),.enable(enable_1[18]),.valid(valid_1[18]),.rdpix(rdpix_1[18]),.addrpix({addrpix_1[82],addrpix_1[18]}));
	pe #(.ADR_WIDTH(2)) pe_1_19 (.state(state_1[79:76]),.ctrlreset(ctrlreset_1[79:76]),.reset(reset_1[79:76]),.enable(enable_1[19]),.valid(valid_1[19]),.rdpix(rdpix_1[19]),.addrpix({addrpix_1[83],addrpix_1[19]}));
	pe #(.ADR_WIDTH(2)) pe_1_20 (.state(state_1[83:80]),.ctrlreset(ctrlreset_1[83:80]),.reset(reset_1[83:80]),.enable(enable_1[20]),.valid(valid_1[20]),.rdpix(rdpix_1[20]),.addrpix({addrpix_1[84],addrpix_1[20]}));
	pe #(.ADR_WIDTH(2)) pe_1_21 (.state(state_1[87:84]),.ctrlreset(ctrlreset_1[87:84]),.reset(reset_1[87:84]),.enable(enable_1[21]),.valid(valid_1[21]),.rdpix(rdpix_1[21]),.addrpix({addrpix_1[85],addrpix_1[21]}));
	pe #(.ADR_WIDTH(2)) pe_1_22 (.state(state_1[91:88]),.ctrlreset(ctrlreset_1[91:88]),.reset(reset_1[91:88]),.enable(enable_1[22]),.valid(valid_1[22]),.rdpix(rdpix_1[22]),.addrpix({addrpix_1[86],addrpix_1[22]}));
	pe #(.ADR_WIDTH(2)) pe_1_23 (.state(state_1[95:92]),.ctrlreset(ctrlreset_1[95:92]),.reset(reset_1[95:92]),.enable(enable_1[23]),.valid(valid_1[23]),.rdpix(rdpix_1[23]),.addrpix({addrpix_1[87],addrpix_1[23]}));
	pe #(.ADR_WIDTH(2)) pe_1_24 (.state(state_1[99:96]),.ctrlreset(ctrlreset_1[99:96]),.reset(reset_1[99:96]),.enable(enable_1[24]),.valid(valid_1[24]),.rdpix(rdpix_1[24]),.addrpix({addrpix_1[88],addrpix_1[24]}));
	pe #(.ADR_WIDTH(2)) pe_1_25 (.state(state_1[103:100]),.ctrlreset(ctrlreset_1[103:100]),.reset(reset_1[103:100]),.enable(enable_1[25]),.valid(valid_1[25]),.rdpix(rdpix_1[25]),.addrpix({addrpix_1[89],addrpix_1[25]}));
	pe #(.ADR_WIDTH(2)) pe_1_26 (.state(state_1[107:104]),.ctrlreset(ctrlreset_1[107:104]),.reset(reset_1[107:104]),.enable(enable_1[26]),.valid(valid_1[26]),.rdpix(rdpix_1[26]),.addrpix({addrpix_1[90],addrpix_1[26]}));
	pe #(.ADR_WIDTH(2)) pe_1_27 (.state(state_1[111:108]),.ctrlreset(ctrlreset_1[111:108]),.reset(reset_1[111:108]),.enable(enable_1[27]),.valid(valid_1[27]),.rdpix(rdpix_1[27]),.addrpix({addrpix_1[91],addrpix_1[27]}));
	pe #(.ADR_WIDTH(2)) pe_1_28 (.state(state_1[115:112]),.ctrlreset(ctrlreset_1[115:112]),.reset(reset_1[115:112]),.enable(enable_1[28]),.valid(valid_1[28]),.rdpix(rdpix_1[28]),.addrpix({addrpix_1[92],addrpix_1[28]}));
	pe #(.ADR_WIDTH(2)) pe_1_29 (.state(state_1[119:116]),.ctrlreset(ctrlreset_1[119:116]),.reset(reset_1[119:116]),.enable(enable_1[29]),.valid(valid_1[29]),.rdpix(rdpix_1[29]),.addrpix({addrpix_1[93],addrpix_1[29]}));
	pe #(.ADR_WIDTH(2)) pe_1_30 (.state(state_1[123:120]),.ctrlreset(ctrlreset_1[123:120]),.reset(reset_1[123:120]),.enable(enable_1[30]),.valid(valid_1[30]),.rdpix(rdpix_1[30]),.addrpix({addrpix_1[94],addrpix_1[30]}));
	pe #(.ADR_WIDTH(2)) pe_1_31 (.state(state_1[127:124]),.ctrlreset(ctrlreset_1[127:124]),.reset(reset_1[127:124]),.enable(enable_1[31]),.valid(valid_1[31]),.rdpix(rdpix_1[31]),.addrpix({addrpix_1[95],addrpix_1[31]}));
	pe #(.ADR_WIDTH(2)) pe_1_32 (.state(state_1[131:128]),.ctrlreset(ctrlreset_1[131:128]),.reset(reset_1[131:128]),.enable(enable_1[32]),.valid(valid_1[32]),.rdpix(rdpix_1[32]),.addrpix({addrpix_1[96],addrpix_1[32]}));
	pe #(.ADR_WIDTH(2)) pe_1_33 (.state(state_1[135:132]),.ctrlreset(ctrlreset_1[135:132]),.reset(reset_1[135:132]),.enable(enable_1[33]),.valid(valid_1[33]),.rdpix(rdpix_1[33]),.addrpix({addrpix_1[97],addrpix_1[33]}));
	pe #(.ADR_WIDTH(2)) pe_1_34 (.state(state_1[139:136]),.ctrlreset(ctrlreset_1[139:136]),.reset(reset_1[139:136]),.enable(enable_1[34]),.valid(valid_1[34]),.rdpix(rdpix_1[34]),.addrpix({addrpix_1[98],addrpix_1[34]}));
	pe #(.ADR_WIDTH(2)) pe_1_35 (.state(state_1[143:140]),.ctrlreset(ctrlreset_1[143:140]),.reset(reset_1[143:140]),.enable(enable_1[35]),.valid(valid_1[35]),.rdpix(rdpix_1[35]),.addrpix({addrpix_1[99],addrpix_1[35]}));
	pe #(.ADR_WIDTH(2)) pe_1_36 (.state(state_1[147:144]),.ctrlreset(ctrlreset_1[147:144]),.reset(reset_1[147:144]),.enable(enable_1[36]),.valid(valid_1[36]),.rdpix(rdpix_1[36]),.addrpix({addrpix_1[100],addrpix_1[36]}));
	pe #(.ADR_WIDTH(2)) pe_1_37 (.state(state_1[151:148]),.ctrlreset(ctrlreset_1[151:148]),.reset(reset_1[151:148]),.enable(enable_1[37]),.valid(valid_1[37]),.rdpix(rdpix_1[37]),.addrpix({addrpix_1[101],addrpix_1[37]}));
	pe #(.ADR_WIDTH(2)) pe_1_38 (.state(state_1[155:152]),.ctrlreset(ctrlreset_1[155:152]),.reset(reset_1[155:152]),.enable(enable_1[38]),.valid(valid_1[38]),.rdpix(rdpix_1[38]),.addrpix({addrpix_1[102],addrpix_1[38]}));
	pe #(.ADR_WIDTH(2)) pe_1_39 (.state(state_1[159:156]),.ctrlreset(ctrlreset_1[159:156]),.reset(reset_1[159:156]),.enable(enable_1[39]),.valid(valid_1[39]),.rdpix(rdpix_1[39]),.addrpix({addrpix_1[103],addrpix_1[39]}));
	pe #(.ADR_WIDTH(2)) pe_1_40 (.state(state_1[163:160]),.ctrlreset(ctrlreset_1[163:160]),.reset(reset_1[163:160]),.enable(enable_1[40]),.valid(valid_1[40]),.rdpix(rdpix_1[40]),.addrpix({addrpix_1[104],addrpix_1[40]}));
	pe #(.ADR_WIDTH(2)) pe_1_41 (.state(state_1[167:164]),.ctrlreset(ctrlreset_1[167:164]),.reset(reset_1[167:164]),.enable(enable_1[41]),.valid(valid_1[41]),.rdpix(rdpix_1[41]),.addrpix({addrpix_1[105],addrpix_1[41]}));
	pe #(.ADR_WIDTH(2)) pe_1_42 (.state(state_1[171:168]),.ctrlreset(ctrlreset_1[171:168]),.reset(reset_1[171:168]),.enable(enable_1[42]),.valid(valid_1[42]),.rdpix(rdpix_1[42]),.addrpix({addrpix_1[106],addrpix_1[42]}));
	pe #(.ADR_WIDTH(2)) pe_1_43 (.state(state_1[175:172]),.ctrlreset(ctrlreset_1[175:172]),.reset(reset_1[175:172]),.enable(enable_1[43]),.valid(valid_1[43]),.rdpix(rdpix_1[43]),.addrpix({addrpix_1[107],addrpix_1[43]}));
	pe #(.ADR_WIDTH(2)) pe_1_44 (.state(state_1[179:176]),.ctrlreset(ctrlreset_1[179:176]),.reset(reset_1[179:176]),.enable(enable_1[44]),.valid(valid_1[44]),.rdpix(rdpix_1[44]),.addrpix({addrpix_1[108],addrpix_1[44]}));
	pe #(.ADR_WIDTH(2)) pe_1_45 (.state(state_1[183:180]),.ctrlreset(ctrlreset_1[183:180]),.reset(reset_1[183:180]),.enable(enable_1[45]),.valid(valid_1[45]),.rdpix(rdpix_1[45]),.addrpix({addrpix_1[109],addrpix_1[45]}));
	pe #(.ADR_WIDTH(2)) pe_1_46 (.state(state_1[187:184]),.ctrlreset(ctrlreset_1[187:184]),.reset(reset_1[187:184]),.enable(enable_1[46]),.valid(valid_1[46]),.rdpix(rdpix_1[46]),.addrpix({addrpix_1[110],addrpix_1[46]}));
	pe #(.ADR_WIDTH(2)) pe_1_47 (.state(state_1[191:188]),.ctrlreset(ctrlreset_1[191:188]),.reset(reset_1[191:188]),.enable(enable_1[47]),.valid(valid_1[47]),.rdpix(rdpix_1[47]),.addrpix({addrpix_1[111],addrpix_1[47]}));
	pe #(.ADR_WIDTH(2)) pe_1_48 (.state(state_1[195:192]),.ctrlreset(ctrlreset_1[195:192]),.reset(reset_1[195:192]),.enable(enable_1[48]),.valid(valid_1[48]),.rdpix(rdpix_1[48]),.addrpix({addrpix_1[112],addrpix_1[48]}));
	pe #(.ADR_WIDTH(2)) pe_1_49 (.state(state_1[199:196]),.ctrlreset(ctrlreset_1[199:196]),.reset(reset_1[199:196]),.enable(enable_1[49]),.valid(valid_1[49]),.rdpix(rdpix_1[49]),.addrpix({addrpix_1[113],addrpix_1[49]}));
	pe #(.ADR_WIDTH(2)) pe_1_50 (.state(state_1[203:200]),.ctrlreset(ctrlreset_1[203:200]),.reset(reset_1[203:200]),.enable(enable_1[50]),.valid(valid_1[50]),.rdpix(rdpix_1[50]),.addrpix({addrpix_1[114],addrpix_1[50]}));
	pe #(.ADR_WIDTH(2)) pe_1_51 (.state(state_1[207:204]),.ctrlreset(ctrlreset_1[207:204]),.reset(reset_1[207:204]),.enable(enable_1[51]),.valid(valid_1[51]),.rdpix(rdpix_1[51]),.addrpix({addrpix_1[115],addrpix_1[51]}));
	pe #(.ADR_WIDTH(2)) pe_1_52 (.state(state_1[211:208]),.ctrlreset(ctrlreset_1[211:208]),.reset(reset_1[211:208]),.enable(enable_1[52]),.valid(valid_1[52]),.rdpix(rdpix_1[52]),.addrpix({addrpix_1[116],addrpix_1[52]}));
	pe #(.ADR_WIDTH(2)) pe_1_53 (.state(state_1[215:212]),.ctrlreset(ctrlreset_1[215:212]),.reset(reset_1[215:212]),.enable(enable_1[53]),.valid(valid_1[53]),.rdpix(rdpix_1[53]),.addrpix({addrpix_1[117],addrpix_1[53]}));
	pe #(.ADR_WIDTH(2)) pe_1_54 (.state(state_1[219:216]),.ctrlreset(ctrlreset_1[219:216]),.reset(reset_1[219:216]),.enable(enable_1[54]),.valid(valid_1[54]),.rdpix(rdpix_1[54]),.addrpix({addrpix_1[118],addrpix_1[54]}));
	pe #(.ADR_WIDTH(2)) pe_1_55 (.state(state_1[223:220]),.ctrlreset(ctrlreset_1[223:220]),.reset(reset_1[223:220]),.enable(enable_1[55]),.valid(valid_1[55]),.rdpix(rdpix_1[55]),.addrpix({addrpix_1[119],addrpix_1[55]}));
	pe #(.ADR_WIDTH(2)) pe_1_56 (.state(state_1[227:224]),.ctrlreset(ctrlreset_1[227:224]),.reset(reset_1[227:224]),.enable(enable_1[56]),.valid(valid_1[56]),.rdpix(rdpix_1[56]),.addrpix({addrpix_1[120],addrpix_1[56]}));
	pe #(.ADR_WIDTH(2)) pe_1_57 (.state(state_1[231:228]),.ctrlreset(ctrlreset_1[231:228]),.reset(reset_1[231:228]),.enable(enable_1[57]),.valid(valid_1[57]),.rdpix(rdpix_1[57]),.addrpix({addrpix_1[121],addrpix_1[57]}));
	pe #(.ADR_WIDTH(2)) pe_1_58 (.state(state_1[235:232]),.ctrlreset(ctrlreset_1[235:232]),.reset(reset_1[235:232]),.enable(enable_1[58]),.valid(valid_1[58]),.rdpix(rdpix_1[58]),.addrpix({addrpix_1[122],addrpix_1[58]}));
	pe #(.ADR_WIDTH(2)) pe_1_59 (.state(state_1[239:236]),.ctrlreset(ctrlreset_1[239:236]),.reset(reset_1[239:236]),.enable(enable_1[59]),.valid(valid_1[59]),.rdpix(rdpix_1[59]),.addrpix({addrpix_1[123],addrpix_1[59]}));
	pe #(.ADR_WIDTH(2)) pe_1_60 (.state(state_1[243:240]),.ctrlreset(ctrlreset_1[243:240]),.reset(reset_1[243:240]),.enable(enable_1[60]),.valid(valid_1[60]),.rdpix(rdpix_1[60]),.addrpix({addrpix_1[124],addrpix_1[60]}));
	pe #(.ADR_WIDTH(2)) pe_1_61 (.state(state_1[247:244]),.ctrlreset(ctrlreset_1[247:244]),.reset(reset_1[247:244]),.enable(enable_1[61]),.valid(valid_1[61]),.rdpix(rdpix_1[61]),.addrpix({addrpix_1[125],addrpix_1[61]}));
	pe #(.ADR_WIDTH(2)) pe_1_62 (.state(state_1[251:248]),.ctrlreset(ctrlreset_1[251:248]),.reset(reset_1[251:248]),.enable(enable_1[62]),.valid(valid_1[62]),.rdpix(rdpix_1[62]),.addrpix({addrpix_1[126],addrpix_1[62]}));
	pe #(.ADR_WIDTH(2)) pe_1_63 (.state(state_1[255:252]),.ctrlreset(ctrlreset_1[255:252]),.reset(reset_1[255:252]),.enable(enable_1[63]),.valid(valid_1[63]),.rdpix(rdpix_1[63]),.addrpix({addrpix_1[127],addrpix_1[63]}));
assign addrpix[3:2] = {|addrpix_1[127:64],|addrpix_1[63:0]};
assign state_1 = valid_0;
assign rdpix_0 = reset_1;
assign enable_0 = ctrlreset_1;
// Level 2
wire [63:0] state_2;
wire [63:0] reset_2;
wire [63:0] ctrlreset_2;
wire [15:0] enable_2;
wire [15:0] rdpix_2;
wire [15:0] valid_2;
wire [31:0] addrpix_2;
	pe #(.ADR_WIDTH(2)) pe_2_0 (.state(state_2[3:0]),.ctrlreset(ctrlreset_2[3:0]),.reset(reset_2[3:0]),.enable(enable_2[0]),.valid(valid_2[0]),.rdpix(rdpix_2[0]),.addrpix({addrpix_2[16],addrpix_2[0]}));
	pe #(.ADR_WIDTH(2)) pe_2_1 (.state(state_2[7:4]),.ctrlreset(ctrlreset_2[7:4]),.reset(reset_2[7:4]),.enable(enable_2[1]),.valid(valid_2[1]),.rdpix(rdpix_2[1]),.addrpix({addrpix_2[17],addrpix_2[1]}));
	pe #(.ADR_WIDTH(2)) pe_2_2 (.state(state_2[11:8]),.ctrlreset(ctrlreset_2[11:8]),.reset(reset_2[11:8]),.enable(enable_2[2]),.valid(valid_2[2]),.rdpix(rdpix_2[2]),.addrpix({addrpix_2[18],addrpix_2[2]}));
	pe #(.ADR_WIDTH(2)) pe_2_3 (.state(state_2[15:12]),.ctrlreset(ctrlreset_2[15:12]),.reset(reset_2[15:12]),.enable(enable_2[3]),.valid(valid_2[3]),.rdpix(rdpix_2[3]),.addrpix({addrpix_2[19],addrpix_2[3]}));
	pe #(.ADR_WIDTH(2)) pe_2_4 (.state(state_2[19:16]),.ctrlreset(ctrlreset_2[19:16]),.reset(reset_2[19:16]),.enable(enable_2[4]),.valid(valid_2[4]),.rdpix(rdpix_2[4]),.addrpix({addrpix_2[20],addrpix_2[4]}));
	pe #(.ADR_WIDTH(2)) pe_2_5 (.state(state_2[23:20]),.ctrlreset(ctrlreset_2[23:20]),.reset(reset_2[23:20]),.enable(enable_2[5]),.valid(valid_2[5]),.rdpix(rdpix_2[5]),.addrpix({addrpix_2[21],addrpix_2[5]}));
	pe #(.ADR_WIDTH(2)) pe_2_6 (.state(state_2[27:24]),.ctrlreset(ctrlreset_2[27:24]),.reset(reset_2[27:24]),.enable(enable_2[6]),.valid(valid_2[6]),.rdpix(rdpix_2[6]),.addrpix({addrpix_2[22],addrpix_2[6]}));
	pe #(.ADR_WIDTH(2)) pe_2_7 (.state(state_2[31:28]),.ctrlreset(ctrlreset_2[31:28]),.reset(reset_2[31:28]),.enable(enable_2[7]),.valid(valid_2[7]),.rdpix(rdpix_2[7]),.addrpix({addrpix_2[23],addrpix_2[7]}));
	pe #(.ADR_WIDTH(2)) pe_2_8 (.state(state_2[35:32]),.ctrlreset(ctrlreset_2[35:32]),.reset(reset_2[35:32]),.enable(enable_2[8]),.valid(valid_2[8]),.rdpix(rdpix_2[8]),.addrpix({addrpix_2[24],addrpix_2[8]}));
	pe #(.ADR_WIDTH(2)) pe_2_9 (.state(state_2[39:36]),.ctrlreset(ctrlreset_2[39:36]),.reset(reset_2[39:36]),.enable(enable_2[9]),.valid(valid_2[9]),.rdpix(rdpix_2[9]),.addrpix({addrpix_2[25],addrpix_2[9]}));
	pe #(.ADR_WIDTH(2)) pe_2_10 (.state(state_2[43:40]),.ctrlreset(ctrlreset_2[43:40]),.reset(reset_2[43:40]),.enable(enable_2[10]),.valid(valid_2[10]),.rdpix(rdpix_2[10]),.addrpix({addrpix_2[26],addrpix_2[10]}));
	pe #(.ADR_WIDTH(2)) pe_2_11 (.state(state_2[47:44]),.ctrlreset(ctrlreset_2[47:44]),.reset(reset_2[47:44]),.enable(enable_2[11]),.valid(valid_2[11]),.rdpix(rdpix_2[11]),.addrpix({addrpix_2[27],addrpix_2[11]}));
	pe #(.ADR_WIDTH(2)) pe_2_12 (.state(state_2[51:48]),.ctrlreset(ctrlreset_2[51:48]),.reset(reset_2[51:48]),.enable(enable_2[12]),.valid(valid_2[12]),.rdpix(rdpix_2[12]),.addrpix({addrpix_2[28],addrpix_2[12]}));
	pe #(.ADR_WIDTH(2)) pe_2_13 (.state(state_2[55:52]),.ctrlreset(ctrlreset_2[55:52]),.reset(reset_2[55:52]),.enable(enable_2[13]),.valid(valid_2[13]),.rdpix(rdpix_2[13]),.addrpix({addrpix_2[29],addrpix_2[13]}));
	pe #(.ADR_WIDTH(2)) pe_2_14 (.state(state_2[59:56]),.ctrlreset(ctrlreset_2[59:56]),.reset(reset_2[59:56]),.enable(enable_2[14]),.valid(valid_2[14]),.rdpix(rdpix_2[14]),.addrpix({addrpix_2[30],addrpix_2[14]}));
	pe #(.ADR_WIDTH(2)) pe_2_15 (.state(state_2[63:60]),.ctrlreset(ctrlreset_2[63:60]),.reset(reset_2[63:60]),.enable(enable_2[15]),.valid(valid_2[15]),.rdpix(rdpix_2[15]),.addrpix({addrpix_2[31],addrpix_2[15]}));
assign addrpix[5:4] = {|addrpix_2[31:16],|addrpix_2[15:0]};
assign state_2 = valid_1;
assign rdpix_1 = reset_2;
assign enable_1 = ctrlreset_2;
// Level 3
wire [15:0] state_3;
wire [15:0] reset_3;
wire [15:0] ctrlreset_3;
wire [3:0] enable_3;
wire [3:0] rdpix_3;
wire [3:0] valid_3;
wire [7:0] addrpix_3;
	pe #(.ADR_WIDTH(2)) pe_3_0 (.state(state_3[3:0]),.ctrlreset(ctrlreset_3[3:0]),.reset(reset_3[3:0]),.enable(enable_3[0]),.valid(valid_3[0]),.rdpix(rdpix_3[0]),.addrpix({addrpix_3[4],addrpix_3[0]}));
	pe #(.ADR_WIDTH(2)) pe_3_1 (.state(state_3[7:4]),.ctrlreset(ctrlreset_3[7:4]),.reset(reset_3[7:4]),.enable(enable_3[1]),.valid(valid_3[1]),.rdpix(rdpix_3[1]),.addrpix({addrpix_3[5],addrpix_3[1]}));
	pe #(.ADR_WIDTH(2)) pe_3_2 (.state(state_3[11:8]),.ctrlreset(ctrlreset_3[11:8]),.reset(reset_3[11:8]),.enable(enable_3[2]),.valid(valid_3[2]),.rdpix(rdpix_3[2]),.addrpix({addrpix_3[6],addrpix_3[2]}));
	pe #(.ADR_WIDTH(2)) pe_3_3 (.state(state_3[15:12]),.ctrlreset(ctrlreset_3[15:12]),.reset(reset_3[15:12]),.enable(enable_3[3]),.valid(valid_3[3]),.rdpix(rdpix_3[3]),.addrpix({addrpix_3[7],addrpix_3[3]}));
assign addrpix[7:6] = {|addrpix_3[7:4],|addrpix_3[3:0]};
assign state_3 = valid_2;
assign rdpix_2 = reset_3;
assign enable_2 = ctrlreset_3;
// Level 4
wire [3:0] state_4;
wire [3:0] reset_4;
wire [3:0] ctrlreset_4;
wire [0:0] enable_4;
wire [0:0] rdpix_4;
wire [0:0] valid_4;
wire [1:0] addrpix_4;
	pe #(.ADR_WIDTH(2)) pe_4_0 (.state(state_4[3:0]),.ctrlreset(ctrlreset_4[3:0]),.reset(reset_4[3:0]),.enable(enable_4[0]),.valid(valid_4[0]),.rdpix(rdpix_4[0]),.addrpix({addrpix_4[1],addrpix_4[0]}));
assign addrpix[9:8] = {|addrpix_4[1:1],|addrpix_4[0:0]};
assign state_4 = valid_3;
assign rdpix_3 = reset_4;
assign enable_3 = ctrlreset_4;
	assign state_0 = state;
	assign reset = reset_0;
	assign rdpix_4 = rdpix;
	assign valid = valid_4;
	assign enable_4 = valid;
endmodule
