
package dut_test_pkg;

`include "dut_test.h"
`include "Packet.sv"
`include "Driver.sv"
`include "Receiver.sv"
`include "Generator.sv"
`include "Scoreboard.sv"
`include "Environment.sv"



endpackage: dut_test_pkg
